// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.10.1.112
// Netlist written on Thu Nov 30 05:38:43 2017
//
// Verilog Description of module vga_leds
//

module vga_leds (CLK50MHZ, hsync, vsync, r, g, b, sram_data, sram_adr, 
            sram_wen, sram_oen, sram_csn) /* synthesis syn_module_defined=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(2[8:16])
    input CLK50MHZ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(3[15:23])
    output hsync;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(5[16:21])
    output vsync;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(6[16:21])
    output [3:0]r;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(9[21:22])
    output [3:0]g;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(10[21:22])
    output [3:0]b;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(11[21:22])
    inout [7:0]sram_data;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(14[20:29])
    output [18:0]sram_adr;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(15[22:30])
    output sram_wen;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(16[16:24])
    output sram_oen;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(17[16:24])
    output sram_csn;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(18[16:24])
    
    wire CLK50MHZ_c /* synthesis is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(3[15:23])
    wire w_clk_video /* synthesis SET_AS_NETWORK=w_clk_video, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(21[6:17])
    wire w_clk_cpu /* synthesis SET_AS_NETWORK=w_clk_cpu, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(22[6:15])
    
    wire GND_net, hsync_c, vsync_c, r_c, r_c_1, r_c_0, g_c, g_c_1, 
        g_c_0, b_c_1, b_c_0, sram_adr_c_18, sram_adr_c_17, sram_adr_c_16, 
        sram_adr_c_15, sram_adr_c_14, sram_adr_c_13, sram_adr_c_12, 
        sram_adr_c_11, sram_adr_c_10, sram_adr_c_9, sram_adr_c_8, sram_adr_c_7, 
        sram_adr_c_6, sram_adr_c_5, sram_adr_c_4, sram_adr_c_3, sram_adr_c_2, 
        sram_adr_c_1, sram_adr_c_0, sram_oen_c, w_locked;
    wire [31:0]counter;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(32[12:19])
    
    wire VCC_net, n23077;
    wire [7:0]sramsram_data_in;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(402[14:30])
    wire [7:0]sramsram_data_out;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(403[14:31])
    wire [2:0]counter_adj_3988;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(428[11:18])
    
    wire reset_n_N_45, n22951, n23112, n22936, n23075, w_clk_cpu_enable_183, 
        n23159, n23099, n23070, n23103, n23156, n23161, n23148, 
        n23175, n23138, n23081, n23083, n23106, n25263, n23127, 
        n23158, n23157, n23072, n23105, n23104, n23150, n23076, 
        n23155, n23147, w_clk_cpu_enable_25, n23124, n42726, n23151, 
        n23060, n23094, n23132, n23183, n23109, n22946;
    wire [4:0]read_idx_0_d;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(470[26:38])
    wire [4:0]read_idx_1_d;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(472[26:38])
    wire [4:0]write_idx_w;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(476[25:36])
    wire [31:0]w_result;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(521[22:30])
    wire [31:0]reg_data_1;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(542[23:33])
    
    wire n23111, n23186, sram_wen_N_3273, n23135, n23092, n23130, 
        n22831, w_clk_cpu_enable_537, n22836, w_clk_cpu_enable_460, 
        n22841, w_clk_cpu_enable_354, n22846, w_clk_cpu_enable_314, 
        n23055, n23071, n23171, n23165, n23064, n22851, n39810, 
        n39809, n23096, n23108, n23153, n39808, w_clk_cpu_enable_23, 
        n22801, n22791, n23139, n23137, n39807, n39806, n39805, 
        n39804, n23174, n39803, n23069, n23101, n23059, n23091, 
        n23163, n23129, n39802, n42732, n42734, n42738, n39801, 
        n39800, n39799, n39798, w_clk_cpu_enable_116, n22956, n39797, 
        n39796, n23078, n23073, w_clk_cpu_enable_279, n23085, n23121, 
        n23173, n23057, w_clk_cpu_enable_323, n23107, n23090, n39773, 
        n23181, n23141, n39772, n23065, n23102, n39771, n39770, 
        n39769, n39768, n39767, n23097, n23134, n23185, n23149, 
        n39766, n39765, n23152, n23140, n39764, n39763, n39762, 
        n39761, n23063, n23084, n23095, n23125, w_clk_cpu_enable_265, 
        n23113, n23160, n23015, n23133, n23123, n23143, w_clk_cpu_enable_107, 
        n23144, n22879, n23074, n23068, n5, n23053, n23087, n23067, 
        n23177, n23167, n5_adj_3986, n22872, n23054, n23061, n23093, 
        n23062, n23052, n39654, n39653, n39652, n39651, n39650, 
        n39649, n39648, n23164, n23145, n22882, n39647, n39646, 
        n39645, n39644, n39643, n39642, n39641, n23162, n23166, 
        n39640, n23142, n23086, n22885, n23146, n23180, n22877, 
        n39625, w_clk_cpu_enable_20, n22874, n22941, n23009, n23082, 
        n23122, w_clk_cpu_enable_576, n23170, n23056, n23089, n22866, 
        n23100, n22926, n23110, w_clk_cpu_enable_188, n41488, n23154, 
        n23172, n23126, n23131, n23176, n41470, n23088, n23182, 
        n23120, n22861, n23079, n23114, n5_adj_3987, w_clk_cpu_enable_137, 
        n23066, n23098, n23080, n22999, n23136, n23178, n22856, 
        n23058, n23115, n23169, n23168, n23128, n23012, n23179;
    
    VHI i6 (.Z(VCC_net));
    BB \u1_1..bidi_cell  (.I(sramsram_data_out[1]), .T(sram_wen_N_3273), 
       .B(sram_data[1]), .O(sramsram_data_in[1])) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=7, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=44 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(408[12] 413[12])
    BB \u1_0..bidi_cell  (.I(sramsram_data_out[0]), .T(sram_wen_N_3273), 
       .B(sram_data[0]), .O(sramsram_data_in[0])) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=7, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=44 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(408[12] 413[12])
    BB \u1_2..bidi_cell  (.I(sramsram_data_out[2]), .T(sram_wen_N_3273), 
       .B(sram_data[2]), .O(sramsram_data_in[2])) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=7, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=44 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(408[12] 413[12])
    BB \u1_3..bidi_cell  (.I(sramsram_data_out[3]), .T(sram_wen_N_3273), 
       .B(sram_data[3]), .O(sramsram_data_in[3])) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=7, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=44 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(408[12] 413[12])
    BB \u1_4..bidi_cell  (.I(sramsram_data_out[4]), .T(sram_wen_N_3273), 
       .B(sram_data[4]), .O(sramsram_data_in[4])) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=7, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=44 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(408[12] 413[12])
    BB \u1_5..bidi_cell  (.I(sramsram_data_out[5]), .T(sram_wen_N_3273), 
       .B(sram_data[5]), .O(sramsram_data_in[5])) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=7, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=44 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(408[12] 413[12])
    BB \u1_6..bidi_cell  (.I(sramsram_data_out[6]), .T(sram_wen_N_3273), 
       .B(sram_data[6]), .O(sramsram_data_in[6])) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=7, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=44 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(408[12] 413[12])
    BB \u1_7..bidi_cell  (.I(sramsram_data_out[7]), .T(sram_wen_N_3273), 
       .B(sram_data[7]), .O(sramsram_data_in[7])) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=7, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=44 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(408[12] 413[12])
    OB sram_adr_pad_16 (.I(sram_adr_c_16), .O(sram_adr[16]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(15[22:30])
    OB sram_adr_pad_17 (.I(sram_adr_c_17), .O(sram_adr[17]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(15[22:30])
    FD1P3AX creset_20477 (.D(n42726), .SP(w_clk_cpu_enable_20), .CK(w_clk_cpu), 
            .Q(n22951));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_20477.GSR = "ENABLED";
    FD1P3AX creset_20381 (.D(n42726), .SP(w_clk_cpu_enable_23), .CK(w_clk_cpu), 
            .Q(n22801));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_20381.GSR = "ENABLED";
    FD1P3AX creset_20449 (.D(n42726), .SP(w_clk_cpu_enable_25), .CK(w_clk_cpu), 
            .Q(n22866));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_20449.GSR = "ENABLED";
    OB sram_adr_pad_18 (.I(sram_adr_c_18), .O(sram_adr[18]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(15[22:30])
    IB CLK50MHZ_pad (.I(CLK50MHZ), .O(CLK50MHZ_c));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(3[15:23])
    OB b_pad_0 (.I(b_c_0), .O(b[0]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(11[21:22])
    OB sram_csn_pad (.I(n41488), .O(sram_csn));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(18[16:24])
    OB b_pad_1 (.I(b_c_1), .O(b[1]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(11[21:22])
    OB sram_oen_pad (.I(sram_oen_c), .O(sram_oen));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(17[16:24])
    OB b_pad_2 (.I(GND_net), .O(b[2]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(11[21:22])
    LUT4 reset_n_I_0_1_lut (.A(w_locked), .Z(reset_n_N_45)) /* synthesis lut_function=(!(A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(431[5:20])
    defparam reset_n_I_0_1_lut.init = 16'h5555;
    PFUMX i37100 (.BLUT(n39652), .ALUT(n39653), .C0(read_idx_0_d[3]), 
          .Z(n39654));
    FD1P3AX creset_20465 (.D(n42726), .SP(w_clk_cpu_enable_107), .CK(w_clk_cpu), 
            .Q(n22936));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_20465.GSR = "ENABLED";
    OB sram_wen_pad (.I(sram_wen_N_3273), .O(sram_wen));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(16[16:24])
    OB b_pad_3 (.I(GND_net), .O(b[3]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(11[21:22])
    FD1P3AX creset_20373 (.D(n42726), .SP(w_clk_cpu_enable_116), .CK(w_clk_cpu), 
            .Q(n22791));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_20373.GSR = "ENABLED";
    OB sram_adr_pad_0 (.I(sram_adr_c_0), .O(sram_adr[0]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(15[22:30])
    OB g_pad_0 (.I(g_c_0), .O(g[0]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(10[21:22])
    OB sram_adr_pad_1 (.I(sram_adr_c_1), .O(sram_adr[1]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(15[22:30])
    OB g_pad_1 (.I(g_c_1), .O(g[1]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(10[21:22])
    FD1P3AX creset_20429 (.D(n42726), .SP(w_clk_cpu_enable_137), .CK(w_clk_cpu), 
            .Q(n22861));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_20429.GSR = "ENABLED";
    OB sram_adr_pad_2 (.I(sram_adr_c_2), .O(sram_adr[2]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(15[22:30])
    OB g_pad_2 (.I(g_c), .O(g[2]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(10[21:22])
    OB sram_adr_pad_3 (.I(sram_adr_c_3), .O(sram_adr[3]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(15[22:30])
    OB g_pad_3 (.I(g_c), .O(g[3]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(10[21:22])
    OB sram_adr_pad_4 (.I(sram_adr_c_4), .O(sram_adr[4]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(15[22:30])
    OB r_pad_0 (.I(r_c_0), .O(r[0]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(9[21:22])
    OB sram_adr_pad_5 (.I(sram_adr_c_5), .O(sram_adr[5]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(15[22:30])
    OB r_pad_1 (.I(r_c_1), .O(r[1]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(9[21:22])
    OB sram_adr_pad_6 (.I(sram_adr_c_6), .O(sram_adr[6]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(15[22:30])
    OB r_pad_2 (.I(r_c), .O(r[2]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(9[21:22])
    OB r_pad_3 (.I(r_c), .O(r[3]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(9[21:22])
    OB sram_adr_pad_7 (.I(sram_adr_c_7), .O(sram_adr[7]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(15[22:30])
    LUT4 i37093_3_lut (.A(n22861), .B(n22866), .C(read_idx_0_d[0]), .Z(n39647)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37093_3_lut.init = 16'hcaca;
    LUT4 i37092_3_lut (.A(n22851), .B(n22856), .C(read_idx_0_d[0]), .Z(n39646)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37092_3_lut.init = 16'hcaca;
    LUT4 i37091_3_lut (.A(n22841), .B(n22846), .C(read_idx_0_d[0]), .Z(n39645)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37091_3_lut.init = 16'hcaca;
    LUT4 i37090_3_lut (.A(n22831), .B(n22836), .C(read_idx_0_d[0]), .Z(n39644)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37090_3_lut.init = 16'hcaca;
    LUT4 i37089_3_lut (.A(n22951), .B(n22956), .C(read_idx_0_d[0]), .Z(n39643)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37089_3_lut.init = 16'hcaca;
    DPR16X4C registers_d01 (.DI0(w_result[28]), .DI1(w_result[29]), .DI2(w_result[30]), 
            .DI3(w_result[31]), .WAD0(n42738), .WAD1(write_idx_w[1]), 
            .WAD2(n42732), .WAD3(n42734), .WCK(w_clk_cpu), .WRE(n23185), 
            .RAD0(read_idx_1_d[0]), .RAD1(read_idx_1_d[1]), .RAD2(read_idx_1_d[2]), 
            .RAD3(read_idx_1_d[3]), .DO0(n23148), .DO1(n23149), .DO2(n23150), 
            .DO3(n23151));
    defparam registers_d01.initval = "0x0000000000000000";
    DPR16X4C registers1 (.DI0(w_result[28]), .DI1(w_result[29]), .DI2(w_result[30]), 
            .DI3(w_result[31]), .WAD0(n42738), .WAD1(write_idx_w[1]), 
            .WAD2(n42732), .WAD3(n42734), .WCK(w_clk_cpu), .WRE(n23185), 
            .RAD0(read_idx_0_d[0]), .RAD1(read_idx_0_d[1]), .RAD2(read_idx_0_d[2]), 
            .RAD3(read_idx_0_d[3]), .DO0(n23080), .DO1(n23081), .DO2(n23082), 
            .DO3(n23083));
    defparam registers1.initval = "0x0000000000000000";
    LUT4 i37088_3_lut (.A(n22941), .B(n22946), .C(read_idx_0_d[0]), .Z(n39642)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37088_3_lut.init = 16'hcaca;
    LUT4 i20526_4_lut (.A(n23009), .B(n39810), .C(n23012), .D(read_idx_1_d[4]), 
         .Z(n23015)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i20526_4_lut.init = 16'hc088;
    LUT4 i37087_3_lut (.A(n22801), .B(n22936), .C(read_idx_0_d[0]), .Z(n39641)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37087_3_lut.init = 16'hcaca;
    FD1P3AX creset_20481 (.D(n42726), .SP(w_clk_cpu_enable_183), .CK(w_clk_cpu), 
            .Q(n22956));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_20481.GSR = "ENABLED";
    LUT4 equal_20514_i2_1_lut (.A(write_idx_w[4]), .Z(n22872)) /* synthesis lut_function=(!(A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam equal_20514_i2_1_lut.init = 16'h5555;
    LUT4 i37086_3_lut (.A(n22791), .B(n22926), .C(read_idx_0_d[0]), .Z(n39640)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37086_3_lut.init = 16'hcaca;
    FD1P3AX creset_20425 (.D(n42726), .SP(w_clk_cpu_enable_188), .CK(w_clk_cpu), 
            .Q(n22856));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_20425.GSR = "ENABLED";
    LUT4 i37219_3_lut (.A(n39770), .B(n39771), .C(write_idx_w[2]), .Z(n39773)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37219_3_lut.init = 16'hcaca;
    LUT4 i37218_3_lut (.A(n39768), .B(n39769), .C(write_idx_w[2]), .Z(n39772)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37218_3_lut.init = 16'hcaca;
    OB sram_adr_pad_8 (.I(sram_adr_c_8), .O(sram_adr[8]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(15[22:30])
    OB sram_adr_pad_9 (.I(sram_adr_c_9), .O(sram_adr[9]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(15[22:30])
    FD1P3AX creset_20421 (.D(n42726), .SP(w_clk_cpu_enable_265), .CK(w_clk_cpu), 
            .Q(n22851));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_20421.GSR = "ENABLED";
    OB sram_adr_pad_10 (.I(sram_adr_c_10), .O(sram_adr[10]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(15[22:30])
    FD1P3AX creset_20457 (.D(n42726), .SP(w_clk_cpu_enable_279), .CK(w_clk_cpu), 
            .Q(n22926));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_20457.GSR = "ENABLED";
    LUT4 equal_20383_i5_2_lut (.A(n42738), .B(write_idx_w[1]), .Z(n5_adj_3987)) /* synthesis lut_function=(A+(B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam equal_20383_i5_2_lut.init = 16'heeee;
    OB sram_adr_pad_11 (.I(sram_adr_c_11), .O(sram_adr[11]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(15[22:30])
    OB sram_adr_pad_12 (.I(sram_adr_c_12), .O(sram_adr[12]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(15[22:30])
    OB vsync_pad (.I(vsync_c), .O(vsync));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(6[16:21])
    OB hsync_pad (.I(hsync_c), .O(hsync));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(5[16:21])
    FD1P3AX creset_20417 (.D(n42726), .SP(w_clk_cpu_enable_314), .CK(w_clk_cpu), 
            .Q(n22846));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_20417.GSR = "ENABLED";
    LUT4 i29723_4_lut (.A(n23122), .B(n23015), .C(n23154), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[2])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29723_4_lut.init = 16'hc088;
    PFUMX i37220 (.BLUT(n39772), .ALUT(n39773), .C0(n42734), .Z(n22999));
    LUT4 i29716_4_lut (.A(n23123), .B(n23015), .C(n23155), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[3])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29716_4_lut.init = 16'hc088;
    FD1P3AX creset_20473 (.D(n42726), .SP(w_clk_cpu_enable_323), .CK(w_clk_cpu), 
            .Q(n22946));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_20473.GSR = "ENABLED";
    LUT4 i29715_4_lut (.A(n23124), .B(n23015), .C(n23156), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[4])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29715_4_lut.init = 16'hc088;
    DPR16X4C n228780 (.DI0(n22872), .DI1(GND_net), .DI2(GND_net), .DI3(GND_net), 
            .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), .WAD2(write_idx_w[2]), 
            .WAD3(n42734), .WCK(w_clk_cpu), .WRE(n22874), .RAD0(read_idx_0_d[0]), 
            .RAD1(read_idx_0_d[1]), .RAD2(read_idx_0_d[2]), .RAD3(read_idx_0_d[3]), 
            .DO0(n22879));
    defparam n228780.initval = "0x0000000000000000";
    FD1P3AX creset_20413 (.D(n42726), .SP(w_clk_cpu_enable_354), .CK(w_clk_cpu), 
            .Q(n22841));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_20413.GSR = "ENABLED";
    DPR16X4C n230110 (.DI0(write_idx_w[4]), .DI1(GND_net), .DI2(GND_net), 
            .DI3(GND_net), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(w_clk_cpu), 
            .WRE(n22877), .RAD0(read_idx_1_d[0]), .RAD1(read_idx_1_d[1]), 
            .RAD2(read_idx_1_d[2]), .RAD3(read_idx_1_d[3]), .DO0(n23012));
    defparam n230110.initval = "0x0000000000000000";
    LUT4 i37249_3_lut (.A(n22861), .B(n22866), .C(read_idx_1_d[0]), .Z(n39803)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37249_3_lut.init = 16'hcaca;
    LUT4 i37248_3_lut (.A(n22851), .B(n22856), .C(read_idx_1_d[0]), .Z(n39802)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37248_3_lut.init = 16'hcaca;
    LUT4 i37247_3_lut (.A(n22841), .B(n22846), .C(read_idx_1_d[0]), .Z(n39801)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37247_3_lut.init = 16'hcaca;
    LUT4 i37246_3_lut (.A(n22831), .B(n22836), .C(read_idx_1_d[0]), .Z(n39800)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37246_3_lut.init = 16'hcaca;
    LUT4 i37245_3_lut (.A(n22951), .B(n22956), .C(read_idx_1_d[0]), .Z(n39799)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37245_3_lut.init = 16'hcaca;
    LUT4 i37244_3_lut (.A(n22941), .B(n22946), .C(read_idx_1_d[0]), .Z(n39798)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37244_3_lut.init = 16'hcaca;
    LUT4 i37243_3_lut (.A(n22801), .B(n22936), .C(read_idx_1_d[0]), .Z(n39797)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37243_3_lut.init = 16'hcaca;
    LUT4 i37242_3_lut (.A(n22791), .B(n22926), .C(read_idx_1_d[0]), .Z(n39796)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37242_3_lut.init = 16'hcaca;
    LUT4 equal_20483_i5_2_lut (.A(n42738), .B(write_idx_w[1]), .Z(n5_adj_3986)) /* synthesis lut_function=((B)+!A) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam equal_20483_i5_2_lut.init = 16'hdddd;
    FD1P3AX creset_20409 (.D(n42726), .SP(w_clk_cpu_enable_460), .CK(w_clk_cpu), 
            .Q(n22836));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_20409.GSR = "ENABLED";
    LUT4 i29706_4_lut (.A(n23125), .B(n23015), .C(n23157), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[5])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29706_4_lut.init = 16'hc088;
    FD1P3AX creset_20405 (.D(n42726), .SP(w_clk_cpu_enable_537), .CK(w_clk_cpu), 
            .Q(n22831));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_20405.GSR = "ENABLED";
    LUT4 i37213_3_lut (.A(n22861), .B(n22866), .C(write_idx_w[0]), .Z(n39767)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37213_3_lut.init = 16'hcaca;
    OB sram_adr_pad_13 (.I(sram_adr_c_13), .O(sram_adr[13]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(15[22:30])
    LUT4 i37212_3_lut (.A(n22851), .B(n22856), .C(write_idx_w[0]), .Z(n39766)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37212_3_lut.init = 16'hcaca;
    FD1P3AX creset_20469 (.D(n42726), .SP(w_clk_cpu_enable_576), .CK(w_clk_cpu), 
            .Q(n22941));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam creset_20469.GSR = "ENABLED";
    LUT4 i37211_3_lut (.A(n22841), .B(n22846), .C(write_idx_w[0]), .Z(n39765)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37211_3_lut.init = 16'hcaca;
    LUT4 i37255_3_lut (.A(n39806), .B(n39807), .C(read_idx_1_d[2]), .Z(n39809)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37255_3_lut.init = 16'hcaca;
    LUT4 i37210_3_lut (.A(n22831), .B(n22836), .C(write_idx_w[0]), .Z(n39764)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37210_3_lut.init = 16'hcaca;
    LUT4 i37209_3_lut (.A(n22951), .B(n22956), .C(write_idx_w[0]), .Z(n39763)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37209_3_lut.init = 16'hcaca;
    LUT4 i37208_3_lut (.A(n22941), .B(n22946), .C(write_idx_w[0]), .Z(n39762)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37208_3_lut.init = 16'hcaca;
    LUT4 i37207_3_lut (.A(n22801), .B(n22936), .C(write_idx_w[0]), .Z(n39761)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37207_3_lut.init = 16'hcaca;
    LUT4 i37071_3_lut (.A(n22791), .B(n22926), .C(write_idx_w[0]), .Z(n39625)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37071_3_lut.init = 16'hcaca;
    LUT4 i37254_3_lut (.A(n39804), .B(n39805), .C(read_idx_1_d[2]), .Z(n39808)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37254_3_lut.init = 16'hcaca;
    LUT4 equal_20407_i5_2_lut (.A(n42738), .B(write_idx_w[1]), .Z(n5)) /* synthesis lut_function=(A+!(B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam equal_20407_i5_2_lut.init = 16'hbbbb;
    LUT4 i1_2_lut_3_lut_4_lut (.A(write_idx_w[3]), .B(n41470), .C(n25263), 
         .D(write_idx_w[2]), .Z(w_clk_cpu_enable_314)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_544 (.A(write_idx_w[3]), .B(n41470), .C(n5), 
         .D(write_idx_w[2]), .Z(w_clk_cpu_enable_354)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_544.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_545 (.A(write_idx_w[3]), .B(n41470), .C(n5_adj_3986), 
         .D(write_idx_w[2]), .Z(w_clk_cpu_enable_460)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_545.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_546 (.A(write_idx_w[3]), .B(n41470), .C(n5_adj_3987), 
         .D(write_idx_w[2]), .Z(w_clk_cpu_enable_537)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_546.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut_adj_547 (.A(write_idx_w[3]), .B(n41470), .C(n25263), 
         .D(write_idx_w[2]), .Z(w_clk_cpu_enable_25)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_547.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_548 (.A(write_idx_w[3]), .B(n41470), .C(n5), 
         .D(write_idx_w[2]), .Z(w_clk_cpu_enable_137)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_548.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_549 (.A(write_idx_w[3]), .B(n41470), .C(n5_adj_3986), 
         .D(write_idx_w[2]), .Z(w_clk_cpu_enable_188)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_549.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut_adj_550 (.A(write_idx_w[3]), .B(n41470), .C(n5_adj_3987), 
         .D(write_idx_w[2]), .Z(w_clk_cpu_enable_265)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_550.init = 16'h0800;
    LUT4 i29179_2_lut (.A(n42738), .B(write_idx_w[1]), .Z(n25263)) /* synthesis lut_function=(A (B)) */ ;
    defparam i29179_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_4_lut_adj_551 (.A(n41470), .B(write_idx_w[3]), .C(n5), 
         .D(write_idx_w[2]), .Z(w_clk_cpu_enable_23)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_551.init = 16'h0002;
    LUT4 i1_2_lut_3_lut_4_lut_adj_552 (.A(n41470), .B(write_idx_w[3]), .C(n25263), 
         .D(write_idx_w[2]), .Z(w_clk_cpu_enable_107)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_552.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_4_lut_adj_553 (.A(n41470), .B(write_idx_w[3]), .C(n5_adj_3987), 
         .D(write_idx_w[2]), .Z(w_clk_cpu_enable_116)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_553.init = 16'h0002;
    LUT4 i1_2_lut_3_lut_4_lut_adj_554 (.A(n41470), .B(write_idx_w[3]), .C(n5_adj_3986), 
         .D(write_idx_w[2]), .Z(w_clk_cpu_enable_279)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_554.init = 16'h0002;
    OB sram_adr_pad_14 (.I(sram_adr_c_14), .O(sram_adr[14]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(15[22:30])
    LUT4 i1_2_lut_3_lut_4_lut_adj_555 (.A(n41470), .B(write_idx_w[3]), .C(n5), 
         .D(write_idx_w[2]), .Z(w_clk_cpu_enable_20)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_555.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_556 (.A(n41470), .B(write_idx_w[3]), .C(n25263), 
         .D(write_idx_w[2]), .Z(w_clk_cpu_enable_183)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_556.init = 16'h2000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_557 (.A(n41470), .B(write_idx_w[3]), .C(n5_adj_3986), 
         .D(write_idx_w[2]), .Z(w_clk_cpu_enable_323)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_557.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_4_lut_adj_558 (.A(n41470), .B(write_idx_w[3]), .C(n5_adj_3987), 
         .D(write_idx_w[2]), .Z(w_clk_cpu_enable_576)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_558.init = 16'h0200;
    LUT4 i37099_3_lut (.A(n39650), .B(n39651), .C(read_idx_0_d[2]), .Z(n39653)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37099_3_lut.init = 16'hcaca;
    PFUMX i37094 (.BLUT(n39640), .ALUT(n39641), .C0(read_idx_0_d[1]), 
          .Z(n39648));
    LUT4 i29724_4_lut (.A(n23121), .B(n23015), .C(n23153), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[1])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29724_4_lut.init = 16'hc088;
    PFUMX i37095 (.BLUT(n39642), .ALUT(n39643), .C0(read_idx_0_d[1]), 
          .Z(n39649));
    PFUMX i37096 (.BLUT(n39644), .ALUT(n39645), .C0(read_idx_0_d[1]), 
          .Z(n39650));
    LUT4 i29705_4_lut (.A(n23126), .B(n23015), .C(n23158), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[6])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29705_4_lut.init = 16'hc088;
    LUT4 i29699_4_lut (.A(n23127), .B(n23015), .C(n23159), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[7])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29699_4_lut.init = 16'hc088;
    PFUMX i37097 (.BLUT(n39646), .ALUT(n39647), .C0(read_idx_0_d[1]), 
          .Z(n39651));
    LUT4 i29698_4_lut (.A(n23128), .B(n23015), .C(n23160), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[8])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29698_4_lut.init = 16'hc088;
    LUT4 i29690_4_lut (.A(n23129), .B(n23015), .C(n23161), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[9])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29690_4_lut.init = 16'hc088;
    LUT4 i29689_4_lut (.A(n23130), .B(n23015), .C(n23162), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[10])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29689_4_lut.init = 16'hc088;
    LUT4 i29682_4_lut (.A(n23131), .B(n23015), .C(n23163), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[11])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29682_4_lut.init = 16'hc088;
    LUT4 i29681_4_lut (.A(n23132), .B(n23015), .C(n23164), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[12])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29681_4_lut.init = 16'hc088;
    LUT4 i29670_4_lut (.A(n23133), .B(n23015), .C(n23165), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[13])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29670_4_lut.init = 16'hc088;
    LUT4 i29669_4_lut (.A(n23134), .B(n23015), .C(n23166), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[14])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29669_4_lut.init = 16'hc088;
    LUT4 i29662_4_lut (.A(n23135), .B(n23015), .C(n23167), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[15])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29662_4_lut.init = 16'hc088;
    LUT4 i29661_4_lut (.A(n23136), .B(n23015), .C(n23168), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[16])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29661_4_lut.init = 16'hc088;
    LUT4 i29649_4_lut (.A(n23137), .B(n23015), .C(n23169), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[17])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29649_4_lut.init = 16'hc088;
    LUT4 i29648_4_lut (.A(n23138), .B(n23015), .C(n23170), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[18])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29648_4_lut.init = 16'hc088;
    LUT4 i29642_4_lut (.A(n23139), .B(n23015), .C(n23171), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[19])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29642_4_lut.init = 16'hc088;
    LUT4 i29641_4_lut (.A(n23140), .B(n23015), .C(n23172), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[20])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29641_4_lut.init = 16'hc088;
    LUT4 i29630_4_lut (.A(n23141), .B(n23015), .C(n23173), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[21])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29630_4_lut.init = 16'hc088;
    LUT4 i29629_4_lut (.A(n23142), .B(n23015), .C(n23174), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[22])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29629_4_lut.init = 16'hc088;
    GSR GSR_INST (.GSR(counter_adj_3988[2]));
    LUT4 i29622_4_lut (.A(n23143), .B(n23015), .C(n23175), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[23])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29622_4_lut.init = 16'hc088;
    LUT4 i29621_4_lut (.A(n23144), .B(n23015), .C(n23176), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[24])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29621_4_lut.init = 16'hc088;
    LUT4 i29614_4_lut (.A(n23145), .B(n23015), .C(n23177), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[25])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29614_4_lut.init = 16'hc088;
    LUT4 i29613_4_lut (.A(n23146), .B(n23015), .C(n23178), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[26])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29613_4_lut.init = 16'hc088;
    VLO i1 (.Z(GND_net));
    TSALL TSALL_INST (.TSALL(GND_net));
    LUT4 i29606_4_lut (.A(n23147), .B(n23015), .C(n23179), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[27])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29606_4_lut.init = 16'hc088;
    LUT4 i29605_4_lut (.A(n23148), .B(n23015), .C(n23180), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[28])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29605_4_lut.init = 16'hc088;
    LUT4 i29593_4_lut (.A(n23149), .B(n23015), .C(n23181), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[29])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29593_4_lut.init = 16'hc088;
    LUT4 i29592_4_lut (.A(n23150), .B(n23015), .C(n23182), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[30])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29592_4_lut.init = 16'hc088;
    LUT4 i29576_4_lut (.A(n23151), .B(n23015), .C(n23183), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[31])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29576_4_lut.init = 16'hc088;
    LUT4 i29711_4_lut (.A(n23120), .B(n23015), .C(n23152), .D(read_idx_1_d[4]), 
         .Z(reg_data_1[0])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i29711_4_lut.init = 16'hc088;
    LUT4 i20446_4_lut (.A(n22879), .B(n39654), .C(n22882), .D(read_idx_0_d[4]), 
         .Z(n22885)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(539[22:31])
    defparam i20446_4_lut.init = 16'hc088;
    DPR16X4C registers_d015 (.DI0(w_result[0]), .DI1(w_result[1]), .DI2(w_result[2]), 
            .DI3(w_result[3]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(w_clk_cpu), 
            .WRE(n23186), .RAD0(read_idx_1_d[0]), .RAD1(read_idx_1_d[1]), 
            .RAD2(read_idx_1_d[2]), .RAD3(read_idx_1_d[3]), .DO0(n23152), 
            .DO1(n23153), .DO2(n23154), .DO3(n23155));
    defparam registers_d015.initval = "0x0000000000000000";
    DPR16X4C registers_d014 (.DI0(w_result[4]), .DI1(w_result[5]), .DI2(w_result[6]), 
            .DI3(w_result[7]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(w_clk_cpu), 
            .WRE(n23186), .RAD0(read_idx_1_d[0]), .RAD1(read_idx_1_d[1]), 
            .RAD2(read_idx_1_d[2]), .RAD3(read_idx_1_d[3]), .DO0(n23156), 
            .DO1(n23157), .DO2(n23158), .DO3(n23159));
    defparam registers_d014.initval = "0x0000000000000000";
    DPR16X4C registers_d013 (.DI0(w_result[8]), .DI1(w_result[9]), .DI2(w_result[10]), 
            .DI3(w_result[11]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(w_clk_cpu), 
            .WRE(n23186), .RAD0(read_idx_1_d[0]), .RAD1(read_idx_1_d[1]), 
            .RAD2(read_idx_1_d[2]), .RAD3(read_idx_1_d[3]), .DO0(n23160), 
            .DO1(n23161), .DO2(n23162), .DO3(n23163));
    defparam registers_d013.initval = "0x0000000000000000";
    DPR16X4C registers_d012 (.DI0(w_result[12]), .DI1(w_result[13]), .DI2(w_result[14]), 
            .DI3(w_result[15]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(w_clk_cpu), 
            .WRE(n23186), .RAD0(read_idx_1_d[0]), .RAD1(read_idx_1_d[1]), 
            .RAD2(read_idx_1_d[2]), .RAD3(read_idx_1_d[3]), .DO0(n23164), 
            .DO1(n23165), .DO2(n23166), .DO3(n23167));
    defparam registers_d012.initval = "0x0000000000000000";
    DPR16X4C registers_d011 (.DI0(w_result[16]), .DI1(w_result[17]), .DI2(w_result[18]), 
            .DI3(w_result[19]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(w_clk_cpu), 
            .WRE(n23186), .RAD0(read_idx_1_d[0]), .RAD1(read_idx_1_d[1]), 
            .RAD2(read_idx_1_d[2]), .RAD3(read_idx_1_d[3]), .DO0(n23168), 
            .DO1(n23169), .DO2(n23170), .DO3(n23171));
    defparam registers_d011.initval = "0x0000000000000000";
    DPR16X4C registers_d010 (.DI0(w_result[20]), .DI1(w_result[21]), .DI2(w_result[22]), 
            .DI3(w_result[23]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(w_clk_cpu), 
            .WRE(n23186), .RAD0(read_idx_1_d[0]), .RAD1(read_idx_1_d[1]), 
            .RAD2(read_idx_1_d[2]), .RAD3(read_idx_1_d[3]), .DO0(n23172), 
            .DO1(n23173), .DO2(n23174), .DO3(n23175));
    defparam registers_d010.initval = "0x0000000000000000";
    DPR16X4C registers_d09 (.DI0(w_result[24]), .DI1(w_result[25]), .DI2(w_result[26]), 
            .DI3(w_result[27]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(w_clk_cpu), 
            .WRE(n23186), .RAD0(read_idx_1_d[0]), .RAD1(read_idx_1_d[1]), 
            .RAD2(read_idx_1_d[2]), .RAD3(read_idx_1_d[3]), .DO0(n23176), 
            .DO1(n23177), .DO2(n23178), .DO3(n23179));
    defparam registers_d09.initval = "0x0000000000000000";
    DPR16X4C registers_d08 (.DI0(w_result[0]), .DI1(w_result[1]), .DI2(w_result[2]), 
            .DI3(w_result[3]), .WAD0(n42738), .WAD1(write_idx_w[1]), .WAD2(n42732), 
            .WAD3(n42734), .WCK(w_clk_cpu), .WRE(n23185), .RAD0(read_idx_1_d[0]), 
            .RAD1(read_idx_1_d[1]), .RAD2(read_idx_1_d[2]), .RAD3(read_idx_1_d[3]), 
            .DO0(n23120), .DO1(n23121), .DO2(n23122), .DO3(n23123));
    defparam registers_d08.initval = "0x0000000000000000";
    DPR16X4C registers_d07 (.DI0(w_result[4]), .DI1(w_result[5]), .DI2(w_result[6]), 
            .DI3(w_result[7]), .WAD0(n42738), .WAD1(write_idx_w[1]), .WAD2(n42732), 
            .WAD3(n42734), .WCK(w_clk_cpu), .WRE(n23185), .RAD0(read_idx_1_d[0]), 
            .RAD1(read_idx_1_d[1]), .RAD2(read_idx_1_d[2]), .RAD3(read_idx_1_d[3]), 
            .DO0(n23124), .DO1(n23125), .DO2(n23126), .DO3(n23127));
    defparam registers_d07.initval = "0x0000000000000000";
    DPR16X4C registers_d06 (.DI0(w_result[8]), .DI1(w_result[9]), .DI2(w_result[10]), 
            .DI3(w_result[11]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(w_clk_cpu), 
            .WRE(n23185), .RAD0(read_idx_1_d[0]), .RAD1(read_idx_1_d[1]), 
            .RAD2(read_idx_1_d[2]), .RAD3(read_idx_1_d[3]), .DO0(n23128), 
            .DO1(n23129), .DO2(n23130), .DO3(n23131));
    defparam registers_d06.initval = "0x0000000000000000";
    DPR16X4C registers_d05 (.DI0(w_result[12]), .DI1(w_result[13]), .DI2(w_result[14]), 
            .DI3(w_result[15]), .WAD0(n42738), .WAD1(write_idx_w[1]), 
            .WAD2(n42732), .WAD3(n42734), .WCK(w_clk_cpu), .WRE(n23185), 
            .RAD0(read_idx_1_d[0]), .RAD1(read_idx_1_d[1]), .RAD2(read_idx_1_d[2]), 
            .RAD3(read_idx_1_d[3]), .DO0(n23132), .DO1(n23133), .DO2(n23134), 
            .DO3(n23135));
    defparam registers_d05.initval = "0x0000000000000000";
    OB sram_adr_pad_15 (.I(sram_adr_c_15), .O(sram_adr[15]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(15[22:30])
    DPR16X4C registers_d04 (.DI0(w_result[16]), .DI1(w_result[17]), .DI2(w_result[18]), 
            .DI3(w_result[19]), .WAD0(n42738), .WAD1(write_idx_w[1]), 
            .WAD2(n42732), .WAD3(n42734), .WCK(w_clk_cpu), .WRE(n23185), 
            .RAD0(read_idx_1_d[0]), .RAD1(read_idx_1_d[1]), .RAD2(read_idx_1_d[2]), 
            .RAD3(read_idx_1_d[3]), .DO0(n23136), .DO1(n23137), .DO2(n23138), 
            .DO3(n23139));
    defparam registers_d04.initval = "0x0000000000000000";
    DPR16X4C registers_d03 (.DI0(w_result[20]), .DI1(w_result[21]), .DI2(w_result[22]), 
            .DI3(w_result[23]), .WAD0(n42738), .WAD1(write_idx_w[1]), 
            .WAD2(n42732), .WAD3(n42734), .WCK(w_clk_cpu), .WRE(n23185), 
            .RAD0(read_idx_1_d[0]), .RAD1(read_idx_1_d[1]), .RAD2(read_idx_1_d[2]), 
            .RAD3(read_idx_1_d[3]), .DO0(n23140), .DO1(n23141), .DO2(n23142), 
            .DO3(n23143));
    defparam registers_d03.initval = "0x0000000000000000";
    DPR16X4C registers_d02 (.DI0(w_result[24]), .DI1(w_result[25]), .DI2(w_result[26]), 
            .DI3(w_result[27]), .WAD0(n42738), .WAD1(write_idx_w[1]), 
            .WAD2(n42732), .WAD3(n42734), .WCK(w_clk_cpu), .WRE(n23185), 
            .RAD0(read_idx_1_d[0]), .RAD1(read_idx_1_d[1]), .RAD2(read_idx_1_d[2]), 
            .RAD3(read_idx_1_d[3]), .DO0(n23144), .DO1(n23145), .DO2(n23146), 
            .DO3(n23147));
    defparam registers_d02.initval = "0x0000000000000000";
    LUT4 i37098_3_lut (.A(n39648), .B(n39649), .C(read_idx_0_d[2]), .Z(n39652)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37098_3_lut.init = 16'hcaca;
    PFUMX i37256 (.BLUT(n39808), .ALUT(n39809), .C0(read_idx_1_d[3]), 
          .Z(n39810));
    DPR16X4C registers15 (.DI0(w_result[0]), .DI1(w_result[1]), .DI2(w_result[2]), 
            .DI3(w_result[3]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(w_clk_cpu), 
            .WRE(n23186), .RAD0(read_idx_0_d[0]), .RAD1(read_idx_0_d[1]), 
            .RAD2(read_idx_0_d[2]), .RAD3(read_idx_0_d[3]), .DO0(n23084), 
            .DO1(n23085), .DO2(n23086), .DO3(n23087));
    defparam registers15.initval = "0x0000000000000000";
    DPR16X4C registers_d00 (.DI0(w_result[28]), .DI1(w_result[29]), .DI2(w_result[30]), 
            .DI3(w_result[31]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(w_clk_cpu), 
            .WRE(n23186), .RAD0(read_idx_1_d[0]), .RAD1(read_idx_1_d[1]), 
            .RAD2(read_idx_1_d[2]), .RAD3(read_idx_1_d[3]), .DO0(n23180), 
            .DO1(n23181), .DO2(n23182), .DO3(n23183));
    defparam registers_d00.initval = "0x0000000000000000";
    DPR16X4C registers14 (.DI0(w_result[4]), .DI1(w_result[5]), .DI2(w_result[6]), 
            .DI3(w_result[7]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(w_clk_cpu), 
            .WRE(n23186), .RAD0(read_idx_0_d[0]), .RAD1(read_idx_0_d[1]), 
            .RAD2(read_idx_0_d[2]), .RAD3(read_idx_0_d[3]), .DO0(n23088), 
            .DO1(n23089), .DO2(n23090), .DO3(n23091));
    defparam registers14.initval = "0x0000000000000000";
    DPR16X4C registers13 (.DI0(w_result[8]), .DI1(w_result[9]), .DI2(w_result[10]), 
            .DI3(w_result[11]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(w_clk_cpu), 
            .WRE(n23186), .RAD0(read_idx_0_d[0]), .RAD1(read_idx_0_d[1]), 
            .RAD2(read_idx_0_d[2]), .RAD3(read_idx_0_d[3]), .DO0(n23092), 
            .DO1(n23093), .DO2(n23094), .DO3(n23095));
    defparam registers13.initval = "0x0000000000000000";
    DPR16X4C registers12 (.DI0(w_result[12]), .DI1(w_result[13]), .DI2(w_result[14]), 
            .DI3(w_result[15]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(w_clk_cpu), 
            .WRE(n23186), .RAD0(read_idx_0_d[0]), .RAD1(read_idx_0_d[1]), 
            .RAD2(read_idx_0_d[2]), .RAD3(read_idx_0_d[3]), .DO0(n23096), 
            .DO1(n23097), .DO2(n23098), .DO3(n23099));
    defparam registers12.initval = "0x0000000000000000";
    DPR16X4C registers11 (.DI0(w_result[16]), .DI1(w_result[17]), .DI2(w_result[18]), 
            .DI3(w_result[19]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(w_clk_cpu), 
            .WRE(n23186), .RAD0(read_idx_0_d[0]), .RAD1(read_idx_0_d[1]), 
            .RAD2(read_idx_0_d[2]), .RAD3(read_idx_0_d[3]), .DO0(n23100), 
            .DO1(n23101), .DO2(n23102), .DO3(n23103));
    defparam registers11.initval = "0x0000000000000000";
    PFUMX i37214 (.BLUT(n39625), .ALUT(n39761), .C0(write_idx_w[1]), .Z(n39768));
    DPR16X4C registers10 (.DI0(w_result[20]), .DI1(w_result[21]), .DI2(w_result[22]), 
            .DI3(w_result[23]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(w_clk_cpu), 
            .WRE(n23186), .RAD0(read_idx_0_d[0]), .RAD1(read_idx_0_d[1]), 
            .RAD2(read_idx_0_d[2]), .RAD3(read_idx_0_d[3]), .DO0(n23104), 
            .DO1(n23105), .DO2(n23106), .DO3(n23107));
    defparam registers10.initval = "0x0000000000000000";
    DPR16X4C registers9 (.DI0(w_result[24]), .DI1(w_result[25]), .DI2(w_result[26]), 
            .DI3(w_result[27]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(w_clk_cpu), 
            .WRE(n23186), .RAD0(read_idx_0_d[0]), .RAD1(read_idx_0_d[1]), 
            .RAD2(read_idx_0_d[2]), .RAD3(read_idx_0_d[3]), .DO0(n23108), 
            .DO1(n23109), .DO2(n23110), .DO3(n23111));
    defparam registers9.initval = "0x0000000000000000";
    DPR16X4C registers8 (.DI0(w_result[0]), .DI1(w_result[1]), .DI2(w_result[2]), 
            .DI3(w_result[3]), .WAD0(n42738), .WAD1(write_idx_w[1]), .WAD2(n42732), 
            .WAD3(n42734), .WCK(w_clk_cpu), .WRE(n23185), .RAD0(read_idx_0_d[0]), 
            .RAD1(read_idx_0_d[1]), .RAD2(read_idx_0_d[2]), .RAD3(read_idx_0_d[3]), 
            .DO0(n23052), .DO1(n23053), .DO2(n23054), .DO3(n23055));
    defparam registers8.initval = "0x0000000000000000";
    DPR16X4C registers7 (.DI0(w_result[4]), .DI1(w_result[5]), .DI2(w_result[6]), 
            .DI3(w_result[7]), .WAD0(n42738), .WAD1(write_idx_w[1]), .WAD2(n42732), 
            .WAD3(n42734), .WCK(w_clk_cpu), .WRE(n23185), .RAD0(read_idx_0_d[0]), 
            .RAD1(read_idx_0_d[1]), .RAD2(read_idx_0_d[2]), .RAD3(read_idx_0_d[3]), 
            .DO0(n23056), .DO1(n23057), .DO2(n23058), .DO3(n23059));
    defparam registers7.initval = "0x0000000000000000";
    DPR16X4C registers6 (.DI0(w_result[8]), .DI1(w_result[9]), .DI2(w_result[10]), 
            .DI3(w_result[11]), .WAD0(n42738), .WAD1(write_idx_w[1]), 
            .WAD2(n42732), .WAD3(n42734), .WCK(w_clk_cpu), .WRE(n23185), 
            .RAD0(read_idx_0_d[0]), .RAD1(read_idx_0_d[1]), .RAD2(read_idx_0_d[2]), 
            .RAD3(read_idx_0_d[3]), .DO0(n23060), .DO1(n23061), .DO2(n23062), 
            .DO3(n23063));
    defparam registers6.initval = "0x0000000000000000";
    DPR16X4C registers5 (.DI0(w_result[12]), .DI1(w_result[13]), .DI2(w_result[14]), 
            .DI3(w_result[15]), .WAD0(n42738), .WAD1(write_idx_w[1]), 
            .WAD2(n42732), .WAD3(n42734), .WCK(w_clk_cpu), .WRE(n23185), 
            .RAD0(read_idx_0_d[0]), .RAD1(read_idx_0_d[1]), .RAD2(read_idx_0_d[2]), 
            .RAD3(read_idx_0_d[3]), .DO0(n23064), .DO1(n23065), .DO2(n23066), 
            .DO3(n23067));
    defparam registers5.initval = "0x0000000000000000";
    PFUMX i37215 (.BLUT(n39762), .ALUT(n39763), .C0(write_idx_w[1]), .Z(n39769));
    DPR16X4C registers4 (.DI0(w_result[16]), .DI1(w_result[17]), .DI2(w_result[18]), 
            .DI3(w_result[19]), .WAD0(n42738), .WAD1(write_idx_w[1]), 
            .WAD2(n42732), .WAD3(n42734), .WCK(w_clk_cpu), .WRE(n23185), 
            .RAD0(read_idx_0_d[0]), .RAD1(read_idx_0_d[1]), .RAD2(read_idx_0_d[2]), 
            .RAD3(read_idx_0_d[3]), .DO0(n23068), .DO1(n23069), .DO2(n23070), 
            .DO3(n23071));
    defparam registers4.initval = "0x0000000000000000";
    DPR16X4C registers3 (.DI0(w_result[20]), .DI1(w_result[21]), .DI2(w_result[22]), 
            .DI3(w_result[23]), .WAD0(n42738), .WAD1(write_idx_w[1]), 
            .WAD2(n42732), .WAD3(n42734), .WCK(w_clk_cpu), .WRE(n23185), 
            .RAD0(read_idx_0_d[0]), .RAD1(read_idx_0_d[1]), .RAD2(read_idx_0_d[2]), 
            .RAD3(read_idx_0_d[3]), .DO0(n23072), .DO1(n23073), .DO2(n23074), 
            .DO3(n23075));
    defparam registers3.initval = "0x0000000000000000";
    DPR16X4C registers2 (.DI0(w_result[24]), .DI1(w_result[25]), .DI2(w_result[26]), 
            .DI3(w_result[27]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(w_clk_cpu), 
            .WRE(n23185), .RAD0(read_idx_0_d[0]), .RAD1(read_idx_0_d[1]), 
            .RAD2(read_idx_0_d[2]), .RAD3(read_idx_0_d[3]), .DO0(n23076), 
            .DO1(n23077), .DO2(n23078), .DO3(n23079));
    defparam registers2.initval = "0x0000000000000000";
    PFUMX i37216 (.BLUT(n39764), .ALUT(n39765), .C0(write_idx_w[1]), .Z(n39770));
    main_pll main_pll_inst (.CLK50MHZ_c(CLK50MHZ_c), .w_clk_video(w_clk_video), 
            .w_clk_cpu(w_clk_cpu), .w_locked(w_locked), .GND_net(GND_net)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(25[10] 30[5])
    PFUMX i37217 (.BLUT(n39766), .ALUT(n39767), .C0(write_idx_w[1]), .Z(n39771));
    display r_3__I_0 (.w_clk_video(w_clk_video), .vsync_c(vsync_c), .hsync_c(hsync_c), 
            .g_c_1(g_c_1), .b_c_1(b_c_1), .g_c_0(g_c_0), .\counter[15] (counter[15]), 
            .\counter[14] (counter[14]), .\counter[13] (counter[13]), .\counter[12] (counter[12]), 
            .\counter[11] (counter[11]), .\counter[10] (counter[10]), .\counter[9] (counter[9]), 
            .\counter[8] (counter[8]), .\counter[7] (counter[7]), .\counter[6] (counter[6]), 
            .\counter[5] (counter[5]), .\counter[4] (counter[4]), .\counter[3] (counter[3]), 
            .\counter[2] (counter[2]), .g_c(g_c), .r_c_1(r_c_1), .r_c(r_c), 
            .\counter[1] (counter[1]), .r_c_0(r_c_0), .b_c_0(b_c_0), .\counter[0] (counter[0]), 
            .reset_n_N_45(reset_n_N_45), .GND_net(GND_net)) /* synthesis syn_module_defined=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(47[9] 58[6])
    DPR16X4C registers0 (.DI0(w_result[28]), .DI1(w_result[29]), .DI2(w_result[30]), 
            .DI3(w_result[31]), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(w_clk_cpu), 
            .WRE(n23186), .RAD0(read_idx_0_d[0]), .RAD1(read_idx_0_d[1]), 
            .RAD2(read_idx_0_d[2]), .RAD3(read_idx_0_d[3]), .DO0(n23112), 
            .DO1(n23113), .DO2(n23114), .DO3(n23115));
    defparam registers0.initval = "0x0000000000000000";
    DPR16X4C n230080 (.DI0(n22872), .DI1(GND_net), .DI2(GND_net), .DI3(GND_net), 
            .WAD0(n42738), .WAD1(write_idx_w[1]), .WAD2(n42732), .WAD3(n42734), 
            .WCK(w_clk_cpu), .WRE(n22874), .RAD0(read_idx_1_d[0]), .RAD1(read_idx_1_d[1]), 
            .RAD2(read_idx_1_d[2]), .RAD3(read_idx_1_d[3]), .DO0(n23009));
    defparam n230080.initval = "0x0000000000000000";
    PFUMX i37250 (.BLUT(n39796), .ALUT(n39797), .C0(read_idx_1_d[1]), 
          .Z(n39804));
    mico_cpu mico_cpu_inst (.\counter[2]_adj_101 (counter_adj_3988[2]), .w_clk_cpu(w_clk_cpu), 
            .reset_n_N_45(reset_n_N_45), .n41488(n41488), .sram_wen_N_3273(sram_wen_N_3273), 
            .n42726(n42726), .sramsram_data_in({sramsram_data_in}), .sram_adr_c_0(sram_adr_c_0), 
            .sramsram_data_out({sramsram_data_out}), .sram_adr_c_18(sram_adr_c_18), 
            .sram_adr_c_17(sram_adr_c_17), .sram_adr_c_16(sram_adr_c_16), 
            .sram_adr_c_15(sram_adr_c_15), .sram_adr_c_14(sram_adr_c_14), 
            .sram_adr_c_13(sram_adr_c_13), .sram_adr_c_12(sram_adr_c_12), 
            .sram_adr_c_11(sram_adr_c_11), .sram_adr_c_10(sram_adr_c_10), 
            .sram_adr_c_9(sram_adr_c_9), .sram_adr_c_8(sram_adr_c_8), .sram_adr_c_7(sram_adr_c_7), 
            .sram_adr_c_6(sram_adr_c_6), .sram_adr_c_5(sram_adr_c_5), .sram_adr_c_4(sram_adr_c_4), 
            .sram_adr_c_3(sram_adr_c_3), .sram_adr_c_2(sram_adr_c_2), .sram_adr_c_1(sram_adr_c_1), 
            .sram_oen_c(sram_oen_c), .\counter[0] (counter[0]), .\counter[1] (counter[1]), 
            .\counter[2] (counter[2]), .\counter[4] (counter[4]), .\counter[5] (counter[5]), 
            .\counter[6] (counter[6]), .\counter[7] (counter[7]), .\counter[8] (counter[8]), 
            .\counter[9] (counter[9]), .\counter[10] (counter[10]), .\counter[11] (counter[11]), 
            .\counter[12] (counter[12]), .\counter[13] (counter[13]), .\counter[14] (counter[14]), 
            .\counter[15] (counter[15]), .\counter[3] (counter[3]), .GND_net(GND_net), 
            .w_result({w_result}), .read_idx_0_d({read_idx_0_d}), .n23059(n23059), 
            .n23091(n23091), .n23058(n23058), .n23090(n23090), .n23067(n23067), 
            .n23099(n23099), .n23068(n23068), .n23100(n23100), .n42734(n42734), 
            .n42738(n42738), .read_idx_1_d({read_idx_1_d}), .n23069(n23069), 
            .n23101(n23101), .n42732(n42732), .n23070(n23070), .n23102(n23102), 
            .n23071(n23071), .n23103(n23103), .n23072(n23072), .n23104(n23104), 
            .n41470(n41470), .write_idx_w({write_idx_w}), .n23185(n23185), 
            .n23186(n23186), .n23073(n23073), .n23105(n23105), .n23074(n23074), 
            .n23106(n23106), .n23075(n23075), .n23107(n23107), .n23076(n23076), 
            .n23108(n23108), .n22885(n22885), .reg_data_1({reg_data_1}), 
            .n23056(n23056), .n23088(n23088), .n23057(n23057), .n23089(n23089), 
            .n22999(n22999), .n22877(n22877), .n22874(n22874), .n23053(n23053), 
            .n23085(n23085), .n23054(n23054), .n23086(n23086), .n23060(n23060), 
            .n23092(n23092), .n23061(n23061), .n23093(n23093), .n23062(n23062), 
            .n23094(n23094), .n23063(n23063), .n23095(n23095), .n23064(n23064), 
            .n23096(n23096), .n23065(n23065), .n23097(n23097), .n23066(n23066), 
            .n23098(n23098), .n23052(n23052), .n23084(n23084), .n23055(n23055), 
            .n23087(n23087), .n23077(n23077), .n23109(n23109), .n23078(n23078), 
            .n23110(n23110), .n23079(n23079), .n23111(n23111), .n23080(n23080), 
            .n23112(n23112), .n23081(n23081), .n23113(n23113), .n23082(n23082), 
            .n23114(n23114), .n23083(n23083), .n23115(n23115), .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(34[10] 44[2])
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    PFUMX i37251 (.BLUT(n39798), .ALUT(n39799), .C0(read_idx_1_d[1]), 
          .Z(n39805));
    DPR16X4C n228810 (.DI0(write_idx_w[4]), .DI1(GND_net), .DI2(GND_net), 
            .DI3(GND_net), .WAD0(write_idx_w[0]), .WAD1(write_idx_w[1]), 
            .WAD2(write_idx_w[2]), .WAD3(write_idx_w[3]), .WCK(w_clk_cpu), 
            .WRE(n22877), .RAD0(read_idx_0_d[0]), .RAD1(read_idx_0_d[1]), 
            .RAD2(read_idx_0_d[2]), .RAD3(read_idx_0_d[3]), .DO0(n22882));
    defparam n228810.initval = "0x0000000000000000";
    PFUMX i37252 (.BLUT(n39800), .ALUT(n39801), .C0(read_idx_1_d[1]), 
          .Z(n39806));
    PFUMX i37253 (.BLUT(n39802), .ALUT(n39803), .C0(read_idx_1_d[1]), 
          .Z(n39807));
    LUT4 m1_lut (.Z(n42726)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module main_pll
//

module main_pll (CLK50MHZ_c, w_clk_video, w_clk_cpu, w_locked, GND_net) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input CLK50MHZ_c;
    output w_clk_video;
    output w_clk_cpu;
    output w_locked;
    input GND_net;
    
    wire CLK50MHZ_c /* synthesis is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(3[15:23])
    wire w_clk_video /* synthesis SET_AS_NETWORK=w_clk_video, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(21[6:17])
    wire w_clk_cpu /* synthesis SET_AS_NETWORK=w_clk_cpu, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(22[6:15])
    
    EHXPLLJ PLLInst_0 (.CLKI(CLK50MHZ_c), .CLKFB(w_clk_video), .PHASESEL0(GND_net), 
            .PHASESEL1(GND_net), .PHASEDIR(GND_net), .PHASESTEP(GND_net), 
            .LOADREG(GND_net), .STDBY(GND_net), .PLLWAKESYNC(GND_net), 
            .RST(GND_net), .RESETC(GND_net), .RESETD(GND_net), .RESETM(GND_net), 
            .ENCLKOP(GND_net), .ENCLKOS(GND_net), .ENCLKOS2(GND_net), 
            .ENCLKOS3(GND_net), .PLLCLK(GND_net), .PLLRST(GND_net), .PLLSTB(GND_net), 
            .PLLWE(GND_net), .PLLDATI0(GND_net), .PLLDATI1(GND_net), .PLLDATI2(GND_net), 
            .PLLDATI3(GND_net), .PLLDATI4(GND_net), .PLLDATI5(GND_net), 
            .PLLDATI6(GND_net), .PLLDATI7(GND_net), .PLLADDR0(GND_net), 
            .PLLADDR1(GND_net), .PLLADDR2(GND_net), .PLLADDR3(GND_net), 
            .PLLADDR4(GND_net), .CLKOP(w_clk_video), .CLKOS(w_clk_cpu), 
            .LOCK(w_locked)) /* synthesis FREQUENCY_PIN_CLKOS="100.000000", FREQUENCY_PIN_CLKOP="75.000000", FREQUENCY_PIN_CLKI="50.000000", ICP_CURRENT="9", LPF_RESISTOR="8", syn_instantiated=1, LSE_LINE_FILE_ID=7, LSE_LCOL=10, LSE_RCOL=5, LSE_LLINE=25, LSE_RLINE=30 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(25[10] 30[5])
    defparam PLLInst_0.CLKI_DIV = 2;
    defparam PLLInst_0.CLKFB_DIV = 3;
    defparam PLLInst_0.CLKOP_DIV = 8;
    defparam PLLInst_0.CLKOS_DIV = 6;
    defparam PLLInst_0.CLKOS2_DIV = 1;
    defparam PLLInst_0.CLKOS3_DIV = 1;
    defparam PLLInst_0.CLKOP_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS_ENABLE = "ENABLED";
    defparam PLLInst_0.CLKOS2_ENABLE = "DISABLED";
    defparam PLLInst_0.CLKOS3_ENABLE = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_A0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_B0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_C0 = "DISABLED";
    defparam PLLInst_0.VCO_BYPASS_D0 = "DISABLED";
    defparam PLLInst_0.CLKOP_CPHASE = 7;
    defparam PLLInst_0.CLKOS_CPHASE = 5;
    defparam PLLInst_0.CLKOS2_CPHASE = 0;
    defparam PLLInst_0.CLKOS3_CPHASE = 0;
    defparam PLLInst_0.CLKOP_FPHASE = 0;
    defparam PLLInst_0.CLKOS_FPHASE = 0;
    defparam PLLInst_0.CLKOS2_FPHASE = 0;
    defparam PLLInst_0.CLKOS3_FPHASE = 0;
    defparam PLLInst_0.FEEDBK_PATH = "CLKOP";
    defparam PLLInst_0.FRACN_ENABLE = "DISABLED";
    defparam PLLInst_0.FRACN_DIV = 0;
    defparam PLLInst_0.CLKOP_TRIM_POL = "RISING";
    defparam PLLInst_0.CLKOP_TRIM_DELAY = 0;
    defparam PLLInst_0.CLKOS_TRIM_POL = "RISING";
    defparam PLLInst_0.CLKOS_TRIM_DELAY = 0;
    defparam PLLInst_0.PLL_USE_WB = "DISABLED";
    defparam PLLInst_0.PREDIVIDER_MUXA1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXB1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXC1 = 0;
    defparam PLLInst_0.PREDIVIDER_MUXD1 = 0;
    defparam PLLInst_0.OUTDIVIDER_MUXA2 = "DIVA";
    defparam PLLInst_0.OUTDIVIDER_MUXB2 = "DIVB";
    defparam PLLInst_0.OUTDIVIDER_MUXC2 = "DIVC";
    defparam PLLInst_0.OUTDIVIDER_MUXD2 = "DIVD";
    defparam PLLInst_0.PLL_LOCK_MODE = 0;
    defparam PLLInst_0.STDBY_ENABLE = "DISABLED";
    defparam PLLInst_0.DPHASE_SOURCE = "DISABLED";
    defparam PLLInst_0.PLLRST_ENA = "DISABLED";
    defparam PLLInst_0.MRST_ENA = "DISABLED";
    defparam PLLInst_0.DCRST_ENA = "DISABLED";
    defparam PLLInst_0.DDRST_ENA = "DISABLED";
    defparam PLLInst_0.INTFB_WAKE = "DISABLED";
    
endmodule
//
// Verilog Description of module display
//

module display (w_clk_video, vsync_c, hsync_c, g_c_1, b_c_1, g_c_0, 
            \counter[15] , \counter[14] , \counter[13] , \counter[12] , 
            \counter[11] , \counter[10] , \counter[9] , \counter[8] , 
            \counter[7] , \counter[6] , \counter[5] , \counter[4] , 
            \counter[3] , \counter[2] , g_c, r_c_1, r_c, \counter[1] , 
            r_c_0, b_c_0, \counter[0] , reset_n_N_45, GND_net) /* synthesis syn_module_defined=1 */ ;
    input w_clk_video;
    output vsync_c;
    output hsync_c;
    output g_c_1;
    output b_c_1;
    output g_c_0;
    input \counter[15] ;
    input \counter[14] ;
    input \counter[13] ;
    input \counter[12] ;
    input \counter[11] ;
    input \counter[10] ;
    input \counter[9] ;
    input \counter[8] ;
    input \counter[7] ;
    input \counter[6] ;
    input \counter[5] ;
    input \counter[4] ;
    input \counter[3] ;
    input \counter[2] ;
    output g_c;
    output r_c_1;
    output r_c;
    input \counter[1] ;
    output r_c_0;
    output b_c_0;
    input \counter[0] ;
    input reset_n_N_45;
    input GND_net;
    
    wire w_clk_video /* synthesis SET_AS_NETWORK=w_clk_video, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(21[6:17])
    wire w_hsync /* synthesis is_clock=1, SET_AS_NETWORK=\r_3__I_0/w_hsync */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(24[6:13])
    wire [6:0]seg7_0;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(127[10:16])
    wire [7:0]seg7_0_6__N_3425;
    
    wire w_vsync, r_vsync_;
    wire [6:0]seg7_1;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(128[10:16])
    wire [7:0]seg7_1_6__N_3432;
    wire [6:0]seg7_2;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(129[10:16])
    wire [7:0]seg7_2_6__N_3439;
    wire [6:0]seg7_3;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(130[10:16])
    wire [7:0]seg7_3_6__N_3446;
    wire [2:0]color_fixed;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(314[10:21])
    wire [2:0]color;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(144[10:15])
    wire [11:0]w_pixel_count;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(27[12:25])
    
    wire n41518, n41448, n4;
    wire [15:0]green_leds_fixed;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(56[25:41])
    
    wire n41519, n202, n41354, n1878, n1431;
    wire [2:0]n1860;
    wire [2:0]n1872;
    
    wire n41355;
    wire [2:0]n1868;
    wire [2:0]n2105;
    
    wire n41487, n4_adj_3976;
    wire [2:0]n1840;
    
    wire vl_seg_line0, vl_seg_line2, n39292;
    wire [2:0]n1168;
    wire [2:0]n2089;
    wire [2:0]n2093;
    
    wire n41358;
    wire [2:0]n2101;
    
    wire n41517, n32565;
    wire [2:0]n2109;
    wire [2:0]color_2__N_3467;
    
    wire n41378, n39417;
    wire [2:0]n1425;
    
    wire n1206;
    wire [2:0]n1421;
    
    wire h_seg_line0, n37517, h_seg_line1, n41449, h_seg_line2, n24, 
        n22, n29675, n40636, n26024, n6, vr_seg_line0;
    wire [2:0]n2113;
    
    wire n41360;
    wire [2:0]n1196;
    wire [2:0]n1188;
    wire [2:0]n1200;
    wire [2:0]color_2__N_3482;
    
    wire n39595, n39788, n36826, n26027, n41379, n39432, n37487, 
        red_leds_fixed_15__N_3476, n39599, vr_seg_line1, n41371, n41350, 
        n41418;
    wire [11:0]w_line_count;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(28[12:24])
    
    wire n41447, n12, n29670, n38917, n39428;
    wire [2:0]n753;
    
    wire n4_adj_3977;
    wire [31:0]n1432;
    wire [2:0]n1864;
    wire [2:0]n1844;
    
    wire vl_seg_line3, n39789, n39790, n41476, n39793, n41489, n41382, 
        n39791, n39792, n39794;
    wire [2:0]n1172;
    
    wire n41381, n41386, n41403;
    wire [2:0]n749;
    
    wire n24_adj_3978, n37473, n565;
    wire [2:0]n1164;
    
    wire n10, n38805;
    wire [2:0]n1836;
    
    wire n24_adj_3979, n41420, n25681, n32490, n534, n24402, n6_adj_3980, 
        n41511, n25680, n32561, n759, n41383, vr_seg_line3;
    wire [2:0]n1848;
    
    wire n41369;
    wire [2:0]n1176;
    
    wire n41404, n38829, n41389, n39164, n16;
    wire [3:0]led_idx;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(78[11:18])
    
    wire n41498, n41521, n14, n32519;
    wire [2:0]n1417;
    
    wire n39524, n31868, n14_adj_3981, n32447, n41415, n41520, n44, 
        n41368, n4_adj_3982, n26020, n32466, n41522;
    wire [2:0]n1192;
    wire [2:0]color_2__N_3470;
    
    wire n41388, n16_adj_3983, n41416;
    wire [2:0]n745;
    
    wire n41617, n41401;
    wire [31:0]color_2__N_3479;
    
    wire n36829, n213, n39782, n39781, n39785, n39784, n39787, 
        n39783, n40635, n4_adj_3984, n39786;
    
    FD1S3AX seg7_0_i0 (.D(seg7_0_6__N_3425[0]), .CK(w_clk_video), .Q(seg7_0[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_0_i0.GSR = "DISABLED";
    FD1S3AX r_vsync_212 (.D(w_vsync), .CK(w_clk_video), .Q(vsync_c)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(59[8] 71[4])
    defparam r_vsync_212.GSR = "DISABLED";
    FD1S3AX r_vsync__213 (.D(vsync_c), .CK(w_clk_video), .Q(r_vsync_)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(59[8] 71[4])
    defparam r_vsync__213.GSR = "DISABLED";
    FD1S3AX seg7_1_i0 (.D(seg7_1_6__N_3432[0]), .CK(w_clk_video), .Q(seg7_1[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_1_i0.GSR = "DISABLED";
    FD1S3AX seg7_2_i0 (.D(seg7_2_6__N_3439[0]), .CK(w_clk_video), .Q(seg7_2[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_2_i0.GSR = "DISABLED";
    FD1S3AX seg7_3_i0 (.D(seg7_3_6__N_3446[0]), .CK(w_clk_video), .Q(seg7_3[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_3_i0.GSR = "DISABLED";
    FD1S3AX color_fixed_i0 (.D(color[0]), .CK(w_clk_video), .Q(color_fixed[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(315[8] 316[21])
    defparam color_fixed_i0.GSR = "DISABLED";
    LUT4 i20253_2_lut_rep_431 (.A(w_pixel_count[0]), .B(w_pixel_count[1]), 
         .Z(n41518)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i20253_2_lut_rep_431.init = 16'heeee;
    LUT4 i20279_2_lut_rep_361_3_lut (.A(w_pixel_count[0]), .B(w_pixel_count[1]), 
         .C(w_pixel_count[2]), .Z(n41448)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i20279_2_lut_rep_361_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut (.A(w_pixel_count[0]), .B(w_pixel_count[1]), .C(w_pixel_count[2]), 
         .Z(n4)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'he0e0;
    LUT4 i33_4_lut (.A(green_leds_fixed[7]), .B(green_leds_fixed[5]), .C(green_leds_fixed[4]), 
         .D(green_leds_fixed[6]), .Z(seg7_1_6__N_3432[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D)))+!A (B (C (D))+!B !(C (D)+!C !(D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(106[2] 123[9])
    defparam i33_4_lut.init = 16'h3ee7;
    FD1S3AX r_hsync_211 (.D(w_hsync), .CK(w_clk_video), .Q(hsync_c)) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(59[8] 71[4])
    defparam r_hsync_211.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_432 (.A(w_pixel_count[6]), .B(w_pixel_count[5]), .Z(n41519)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_432.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_517 (.A(w_pixel_count[6]), .B(w_pixel_count[5]), 
         .C(w_pixel_count[7]), .Z(n202)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;
    defparam i1_2_lut_3_lut_adj_517.init = 16'hf8f8;
    LUT4 green_leds_fixed_4__bdd_4_lut (.A(green_leds_fixed[4]), .B(green_leds_fixed[7]), 
         .C(green_leds_fixed[6]), .D(green_leds_fixed[5]), .Z(seg7_1_6__N_3432[4])) /* synthesis lut_function=(A (B (C+(D)))+!A (B+((D)+!C))) */ ;
    defparam green_leds_fixed_4__bdd_4_lut.init = 16'hddc5;
    LUT4 green_leds_fixed_13__bdd_4_lut_38457 (.A(green_leds_fixed[13]), .B(green_leds_fixed[12]), 
         .C(green_leds_fixed[15]), .D(green_leds_fixed[14]), .Z(seg7_3_6__N_3446[5])) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A !(B (C (D)+!C !(D)))) */ ;
    defparam green_leds_fixed_13__bdd_4_lut_38457.init = 16'hb7f1;
    FD1S3AX seg7_1_i6 (.D(seg7_1_6__N_3432[6]), .CK(w_clk_video), .Q(seg7_1[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_1_i6.GSR = "DISABLED";
    LUT4 i37630_3_lut_4_lut (.A(n41354), .B(n1878), .C(n1431), .D(n1860[0]), 
         .Z(n1872[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(311[3:11])
    defparam i37630_3_lut_4_lut.init = 16'h8f80;
    FD1S3AX seg7_1_i5 (.D(seg7_1_6__N_3432[5]), .CK(w_clk_video), .Q(seg7_1[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_1_i5.GSR = "DISABLED";
    LUT4 i37635_3_lut_4_lut_4_lut (.A(n41355), .B(n1868[0]), .C(n1872[0]), 
         .D(n1431), .Z(n2105[0])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(288[2] 311[11])
    defparam i37635_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 mux_9_Mux_2_i15_4_lut (.A(green_leds_fixed[6]), .B(green_leds_fixed[4]), 
         .C(green_leds_fixed[7]), .D(green_leds_fixed[5]), .Z(seg7_1_6__N_3432[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A !(B+(C+!(D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(106[2] 123[9])
    defparam mux_9_Mux_2_i15_4_lut.init = 16'h5edf;
    FD1S3AX seg7_1_i4 (.D(seg7_1_6__N_3432[4]), .CK(w_clk_video), .Q(seg7_1[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_1_i4.GSR = "DISABLED";
    FD1S3AX seg7_1_i3 (.D(seg7_1_6__N_3432[3]), .CK(w_clk_video), .Q(seg7_1[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_1_i3.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_3_lut (.A(color_fixed[0]), .B(color_fixed[2]), .C(color_fixed[1]), 
         .Z(g_c_1)) /* synthesis lut_function=(A (B+!(C))+!A (C)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(315[8] 316[21])
    defparam i1_2_lut_3_lut_3_lut.init = 16'hdada;
    FD1S3AX seg7_1_i2 (.D(seg7_1_6__N_3432[2]), .CK(w_clk_video), .Q(seg7_1[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_1_i2.GSR = "DISABLED";
    LUT4 mux_175_i1_3_lut_4_lut (.A(n41487), .B(n4_adj_3976), .C(seg7_1[4]), 
         .D(seg7_2[4]), .Z(n1840[0])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_175_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 i38090_2_lut_3_lut_4_lut (.A(n41487), .B(n4_adj_3976), .C(vl_seg_line0), 
         .D(vl_seg_line2), .Z(n39292)) /* synthesis lut_function=(A (C+(D))+!A (B+(C+(D)))) */ ;
    defparam i38090_2_lut_3_lut_4_lut.init = 16'hfff4;
    FD1S3AX seg7_1_i1 (.D(seg7_1_6__N_3432[1]), .CK(w_clk_video), .Q(seg7_1[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_1_i1.GSR = "DISABLED";
    FD1S3AX seg7_0_i6 (.D(seg7_0_6__N_3425[6]), .CK(w_clk_video), .Q(seg7_0[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_0_i6.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut_adj_518 (.A(color_fixed[0]), .B(color_fixed[2]), 
         .C(color_fixed[1]), .Z(b_c_1)) /* synthesis lut_function=(A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(315[8] 316[21])
    defparam i1_2_lut_3_lut_adj_518.init = 16'h8080;
    LUT4 mux_133_i1_3_lut_4_lut (.A(n41487), .B(n4_adj_3976), .C(seg7_1[5]), 
         .D(seg7_2[5]), .Z(n1168[0])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_133_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_4_lut_3_lut (.A(color_fixed[0]), .B(color_fixed[2]), .C(color_fixed[1]), 
         .Z(g_c_0)) /* synthesis lut_function=(A (B+!(C))+!A ((C)+!B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(315[8] 316[21])
    defparam i1_4_lut_3_lut.init = 16'hdbdb;
    LUT4 i29174_2_lut_4_lut (.A(n2089[1]), .B(n2093[1]), .C(n41358), .D(n1878), 
         .Z(n2101[1])) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i29174_2_lut_4_lut.init = 16'hca00;
    FD1S3AX seg7_0_i5 (.D(seg7_0_6__N_3425[5]), .CK(w_clk_video), .Q(seg7_0[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_0_i5.GSR = "DISABLED";
    LUT4 i29981_4_lut (.A(n41517), .B(n4), .C(w_pixel_count[4]), .D(w_pixel_count[3]), 
         .Z(n32565)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i29981_4_lut.init = 16'hfaea;
    FD1S3AX seg7_0_i4 (.D(seg7_0_6__N_3425[4]), .CK(w_clk_video), .Q(seg7_0[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_0_i4.GSR = "DISABLED";
    LUT4 color_2__I_0_i2_4_lut (.A(n2109[1]), .B(color_2__N_3467[1]), .C(n41378), 
         .D(n39417), .Z(color[1])) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(155[2] 311[11])
    defparam color_2__I_0_i2_4_lut.init = 16'hcacc;
    LUT4 mux_201_i2_3_lut (.A(n2105[1]), .B(n1425[1]), .C(n1206), .Z(n2109[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(248[2] 311[11])
    defparam mux_201_i2_3_lut.init = 16'hcaca;
    LUT4 mux_156_i2_3_lut (.A(n1421[1]), .B(seg7_0[6]), .C(h_seg_line0), 
         .Z(n1425[1])) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(230[3] 245[12])
    defparam mux_156_i2_3_lut.init = 16'h3a3a;
    LUT4 mux_155_i2_3_lut (.A(n37517), .B(seg7_1[6]), .C(h_seg_line1), 
         .Z(n1421[1])) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(233[3] 245[12])
    defparam mux_155_i2_3_lut.init = 16'h3a3a;
    LUT4 i42_4_lut (.A(n41449), .B(seg7_2[6]), .C(h_seg_line2), .D(n24), 
         .Z(n37517)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(236[3] 245[12])
    defparam i42_4_lut.init = 16'h3a30;
    LUT4 i43_4_lut (.A(n22), .B(n29675), .C(w_pixel_count[7]), .D(seg7_3[6]), 
         .Z(n24)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(236[3] 245[12])
    defparam i43_4_lut.init = 16'h0aca;
    LUT4 mux_11_Mux_2_i15_4_lut (.A(green_leds_fixed[14]), .B(green_leds_fixed[12]), 
         .C(green_leds_fixed[15]), .D(green_leds_fixed[13]), .Z(seg7_3_6__N_3446[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A !(B+(C+!(D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(106[2] 123[9])
    defparam mux_11_Mux_2_i15_4_lut.init = 16'h5edf;
    LUT4 i29163_4_lut (.A(n40636), .B(n26024), .C(n6), .D(vr_seg_line0), 
         .Z(n2113[2])) /* synthesis lut_function=(A (B)+!A (B (C+(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(225[2] 311[11])
    defparam i29163_4_lut.init = 16'hccc8;
    LUT4 mux_10_Mux_2_i15_4_lut (.A(green_leds_fixed[10]), .B(green_leds_fixed[8]), 
         .C(green_leds_fixed[11]), .D(green_leds_fixed[9]), .Z(seg7_2_6__N_3439[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A !(B+(C+!(D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(106[2] 123[9])
    defparam mux_10_Mux_2_i15_4_lut.init = 16'h5edf;
    LUT4 i37632_3_lut_4_lut (.A(vr_seg_line0), .B(n41360), .C(n1196[0]), 
         .D(n1188[0]), .Z(n1200[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(189[3] 222[12])
    defparam i37632_3_lut_4_lut.init = 16'hf1e0;
    L6MUX21 i36509 (.D0(n2109[0]), .D1(color_2__N_3482[0]), .SD(n39595), 
            .Z(color[0]));
    LUT4 i37234_3_lut_3_lut (.A(w_pixel_count[5]), .B(green_leds_fixed[7]), 
         .C(green_leds_fixed[6]), .Z(n39788)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(78[37:70])
    defparam i37234_3_lut_3_lut.init = 16'he4e4;
    FD1S3AX seg7_0_i3 (.D(seg7_0_6__N_3425[3]), .CK(w_clk_video), .Q(seg7_0[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_0_i3.GSR = "DISABLED";
    PFUMX mux_201_i1 (.BLUT(n2105[0]), .ALUT(n1425[0]), .C0(n1206), .Z(n2109[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;
    FD1S3AX seg7_0_i2 (.D(seg7_0_6__N_3425[2]), .CK(w_clk_video), .Q(seg7_0[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_0_i2.GSR = "DISABLED";
    PFUMX mux_203_i3 (.BLUT(n2113[2]), .ALUT(n36826), .C0(n26027), .Z(color_2__N_3482[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;
    FD1S3AX seg7_0_i1 (.D(seg7_0_6__N_3425[1]), .CK(w_clk_video), .Q(seg7_0[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_0_i1.GSR = "DISABLED";
    LUT4 i38073_2_lut_rep_271 (.A(h_seg_line0), .B(h_seg_line1), .Z(n41358)) /* synthesis lut_function=(A+(B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(167[3] 182[12])
    defparam i38073_2_lut_rep_271.init = 16'heeee;
    LUT4 i38037_3_lut_3_lut_4_lut (.A(h_seg_line0), .B(h_seg_line1), .C(n41378), 
         .D(n41379), .Z(n39432)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(167[3] 182[12])
    defparam i38037_3_lut_3_lut_4_lut.init = 16'hf0f1;
    LUT4 i37593_3_lut_rep_267_4_lut (.A(h_seg_line0), .B(h_seg_line1), .C(n2093[0]), 
         .D(n37487), .Z(n41354)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(167[3] 182[12])
    defparam i37593_3_lut_rep_267_4_lut.init = 16'hf1e0;
    FD1P3AX green_leds_fixed_i0_i15 (.D(\counter[15] ), .SP(red_leds_fixed_15__N_3476), 
            .CK(w_clk_video), .Q(green_leds_fixed[15])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(59[8] 71[4])
    defparam green_leds_fixed_i0_i15.GSR = "DISABLED";
    FD1P3AX green_leds_fixed_i0_i14 (.D(\counter[14] ), .SP(red_leds_fixed_15__N_3476), 
            .CK(w_clk_video), .Q(green_leds_fixed[14])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(59[8] 71[4])
    defparam green_leds_fixed_i0_i14.GSR = "DISABLED";
    FD1P3AX green_leds_fixed_i0_i13 (.D(\counter[13] ), .SP(red_leds_fixed_15__N_3476), 
            .CK(w_clk_video), .Q(green_leds_fixed[13])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(59[8] 71[4])
    defparam green_leds_fixed_i0_i13.GSR = "DISABLED";
    FD1P3AX green_leds_fixed_i0_i12 (.D(\counter[12] ), .SP(red_leds_fixed_15__N_3476), 
            .CK(w_clk_video), .Q(green_leds_fixed[12])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(59[8] 71[4])
    defparam green_leds_fixed_i0_i12.GSR = "DISABLED";
    FD1P3AX green_leds_fixed_i0_i11 (.D(\counter[11] ), .SP(red_leds_fixed_15__N_3476), 
            .CK(w_clk_video), .Q(green_leds_fixed[11])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(59[8] 71[4])
    defparam green_leds_fixed_i0_i11.GSR = "DISABLED";
    FD1P3AX green_leds_fixed_i0_i10 (.D(\counter[10] ), .SP(red_leds_fixed_15__N_3476), 
            .CK(w_clk_video), .Q(green_leds_fixed[10])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(59[8] 71[4])
    defparam green_leds_fixed_i0_i10.GSR = "DISABLED";
    PFUMX mux_203_i1 (.BLUT(n1200[0]), .ALUT(n2113[0]), .C0(n39599), .Z(color_2__N_3482[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;
    FD1P3AX green_leds_fixed_i0_i9 (.D(\counter[9] ), .SP(red_leds_fixed_15__N_3476), 
            .CK(w_clk_video), .Q(green_leds_fixed[9])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(59[8] 71[4])
    defparam green_leds_fixed_i0_i9.GSR = "DISABLED";
    FD1P3AX green_leds_fixed_i0_i8 (.D(\counter[8] ), .SP(red_leds_fixed_15__N_3476), 
            .CK(w_clk_video), .Q(green_leds_fixed[8])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(59[8] 71[4])
    defparam green_leds_fixed_i0_i8.GSR = "DISABLED";
    FD1P3AX green_leds_fixed_i0_i7 (.D(\counter[7] ), .SP(red_leds_fixed_15__N_3476), 
            .CK(w_clk_video), .Q(green_leds_fixed[7])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(59[8] 71[4])
    defparam green_leds_fixed_i0_i7.GSR = "DISABLED";
    FD1P3AX green_leds_fixed_i0_i6 (.D(\counter[6] ), .SP(red_leds_fixed_15__N_3476), 
            .CK(w_clk_video), .Q(green_leds_fixed[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(59[8] 71[4])
    defparam green_leds_fixed_i0_i6.GSR = "DISABLED";
    FD1P3AX green_leds_fixed_i0_i5 (.D(\counter[5] ), .SP(red_leds_fixed_15__N_3476), 
            .CK(w_clk_video), .Q(green_leds_fixed[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(59[8] 71[4])
    defparam green_leds_fixed_i0_i5.GSR = "DISABLED";
    FD1P3AX green_leds_fixed_i0_i4 (.D(\counter[4] ), .SP(red_leds_fixed_15__N_3476), 
            .CK(w_clk_video), .Q(green_leds_fixed[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(59[8] 71[4])
    defparam green_leds_fixed_i0_i4.GSR = "DISABLED";
    LUT4 i37834_2_lut_rep_268_3_lut (.A(vr_seg_line1), .B(n41371), .C(vr_seg_line0), 
         .Z(n41355)) /* synthesis lut_function=(A+(B+(C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(189[3] 222[12])
    defparam i37834_2_lut_rep_268_3_lut.init = 16'hfefe;
    LUT4 i37843_2_lut_rep_263_2_lut_3_lut_4_lut (.A(vr_seg_line1), .B(n41371), 
         .C(n1431), .D(vr_seg_line0), .Z(n41350)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+!(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(189[3] 222[12])
    defparam i37843_2_lut_rep_263_2_lut_3_lut_4_lut.init = 16'hf0f1;
    LUT4 i1_2_lut_rep_331_3_lut_4_lut (.A(w_pixel_count[4]), .B(w_pixel_count[3]), 
         .C(w_pixel_count[2]), .D(n41518), .Z(n41418)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i1_2_lut_rep_331_3_lut_4_lut.init = 16'h8880;
    FD1P3AX green_leds_fixed_i0_i3 (.D(\counter[3] ), .SP(red_leds_fixed_15__N_3476), 
            .CK(w_clk_video), .Q(green_leds_fixed[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(59[8] 71[4])
    defparam green_leds_fixed_i0_i3.GSR = "DISABLED";
    FD1P3AX green_leds_fixed_i0_i2 (.D(\counter[2] ), .SP(red_leds_fixed_15__N_3476), 
            .CK(w_clk_video), .Q(green_leds_fixed[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(59[8] 71[4])
    defparam green_leds_fixed_i0_i2.GSR = "DISABLED";
    LUT4 i1_2_lut (.A(color_fixed[1]), .B(color_fixed[0]), .Z(g_c)) /* synthesis lut_function=(!(A+!(B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(315[8] 316[21])
    defparam i1_2_lut.init = 16'h4444;
    LUT4 i20339_2_lut_4_lut (.A(w_line_count[3]), .B(w_line_count[4]), .C(n41447), 
         .D(w_line_count[5]), .Z(n12)) /* synthesis lut_function=(A (B+(D))+!A (B (C+(D))+!B (D))) */ ;
    defparam i20339_2_lut_4_lut.init = 16'hffc8;
    LUT4 i1_3_lut_4_lut (.A(w_pixel_count[3]), .B(n41448), .C(w_pixel_count[4]), 
         .D(w_pixel_count[5]), .Z(n29670)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C (D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hfe00;
    LUT4 i1_4_lut_4_lut (.A(w_pixel_count[3]), .B(n41448), .C(w_pixel_count[4]), 
         .D(w_pixel_count[5]), .Z(n22)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (D)+!B (C (D))))) */ ;
    defparam i1_4_lut_4_lut.init = 16'h5e00;
    LUT4 i1_3_lut (.A(color_fixed[1]), .B(color_fixed[2]), .C(color_fixed[0]), 
         .Z(r_c_1)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(314[10:21])
    defparam i1_3_lut.init = 16'hecec;
    LUT4 i2_3_lut_4_lut (.A(w_pixel_count[7]), .B(n41449), .C(n38917), 
         .D(w_pixel_count[6]), .Z(h_seg_line2)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_3_lut_adj_519 (.A(color_fixed[0]), .B(color_fixed[2]), .C(color_fixed[1]), 
         .Z(r_c)) /* synthesis lut_function=(!((B (C)+!B !(C))+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(315[8] 316[21])
    defparam i1_3_lut_adj_519.init = 16'h2828;
    FD1P3AX green_leds_fixed_i0_i1 (.D(\counter[1] ), .SP(red_leds_fixed_15__N_3476), 
            .CK(w_clk_video), .Q(green_leds_fixed[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(59[8] 71[4])
    defparam green_leds_fixed_i0_i1.GSR = "DISABLED";
    L6MUX21 mux_200_i2 (.D0(n1868[1]), .D1(n1872[1]), .SD(n41350), .Z(n2105[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;
    L6MUX21 color_2__I_173_i2 (.D0(n1200[1]), .D1(color_2__N_3482[1]), .SD(n39428), 
            .Z(color_2__N_3467[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;
    LUT4 green_leds_fixed_12__bdd_4_lut (.A(green_leds_fixed[12]), .B(green_leds_fixed[15]), 
         .C(green_leds_fixed[13]), .D(green_leds_fixed[14]), .Z(seg7_3_6__N_3446[0])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+(D)))+!A (B+(C+!(D)))) */ ;
    defparam green_leds_fixed_12__bdd_4_lut.init = 16'hf67d;
    PFUMX mux_141_i2 (.BLUT(n1188[1]), .ALUT(n1196[1]), .C0(n41355), .Z(n1200[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;
    PFUMX mux_183_i2 (.BLUT(n1860[1]), .ALUT(n2101[1]), .C0(n1431), .Z(n1872[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;
    PFUMX mux_203_i2 (.BLUT(n753[1]), .ALUT(n2113[1]), .C0(n39432), .Z(color_2__N_3482[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;
    LUT4 w_pixel_count_6__bdd_4_lut_38833 (.A(w_pixel_count[6]), .B(n41418), 
         .C(w_pixel_count[7]), .D(w_pixel_count[5]), .Z(n4_adj_3977)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam w_pixel_count_6__bdd_4_lut_38833.init = 16'h0008;
    LUT4 i53_1_lut (.A(seg7_0[2]), .Z(n1432[1])) /* synthesis lut_function=(!(A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(250[12:29])
    defparam i53_1_lut.init = 16'h5555;
    LUT4 mux_181_i2_3_lut (.A(seg7_2[2]), .B(seg7_1[2]), .C(vr_seg_line1), 
         .Z(n1864[1])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(258[3] 285[12])
    defparam mux_181_i2_3_lut.init = 16'h3535;
    LUT4 mux_176_i2_3_lut (.A(seg7_1[4]), .B(seg7_0[4]), .C(vl_seg_line0), 
         .Z(n1844[1])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(273[3] 285[12])
    defparam mux_176_i2_3_lut.init = 16'h3535;
    LUT4 mux_175_i2_4_lut (.A(seg7_3[4]), .B(seg7_2[4]), .C(vl_seg_line2), 
         .D(vl_seg_line3), .Z(n1840[1])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(276[3] 285[12])
    defparam mux_175_i2_4_lut.init = 16'h3530;
    LUT4 green_leds_fixed_12__bdd_4_lut_38522 (.A(green_leds_fixed[12]), .B(green_leds_fixed[15]), 
         .C(green_leds_fixed[14]), .D(green_leds_fixed[13]), .Z(seg7_3_6__N_3446[4])) /* synthesis lut_function=(A (B (C+(D)))+!A (B+((D)+!C))) */ ;
    defparam green_leds_fixed_12__bdd_4_lut_38522.init = 16'hddc5;
    LUT4 w_pixel_count_3__bdd_4_lut (.A(w_pixel_count[3]), .B(w_pixel_count[5]), 
         .C(w_pixel_count[4]), .D(n41448), .Z(n38917)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C+(D))))) */ ;
    defparam w_pixel_count_3__bdd_4_lut.init = 16'h4c48;
    L6MUX21 i37239 (.D0(n39789), .D1(n39790), .SD(n41476), .Z(n39793));
    LUT4 i20219_2_lut_rep_295_3_lut_4_lut (.A(n41448), .B(n41489), .C(w_pixel_count[6]), 
         .D(w_pixel_count[5]), .Z(n41382)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i20219_2_lut_rep_295_3_lut_4_lut.init = 16'hfff8;
    L6MUX21 i37240 (.D0(n39791), .D1(n39792), .SD(n41476), .Z(n39794));
    LUT4 mux_134_i2_3_lut (.A(seg7_1[5]), .B(seg7_0[5]), .C(vl_seg_line0), 
         .Z(n1172[1])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(210[3] 222[12])
    defparam mux_134_i2_3_lut.init = 16'h3535;
    LUT4 mux_133_i2_4_lut (.A(seg7_3[5]), .B(seg7_2[5]), .C(vl_seg_line2), 
         .D(vl_seg_line3), .Z(n1168[1])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(213[3] 222[12])
    defparam mux_133_i2_4_lut.init = 16'h3530;
    LUT4 i20268_2_lut_rep_294_3_lut_4_lut (.A(n41448), .B(n41489), .C(w_pixel_count[6]), 
         .D(w_pixel_count[5]), .Z(n41381)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i20268_2_lut_rep_294_3_lut_4_lut.init = 16'hf080;
    LUT4 green_leds_fixed_8__bdd_4_lut_38527 (.A(green_leds_fixed[8]), .B(green_leds_fixed[11]), 
         .C(green_leds_fixed[10]), .D(green_leds_fixed[9]), .Z(seg7_2_6__N_3439[4])) /* synthesis lut_function=(A (B (C+(D)))+!A (B+((D)+!C))) */ ;
    defparam green_leds_fixed_8__bdd_4_lut_38527.init = 16'hddc5;
    LUT4 i20285_2_lut_rep_299_3_lut_4_lut (.A(n41448), .B(n41489), .C(w_pixel_count[6]), 
         .D(w_pixel_count[5]), .Z(n41386)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20285_2_lut_rep_299_3_lut_4_lut.init = 16'h8000;
    LUT4 vr_seg_line2_I_0_3_lut_rep_284_4_lut (.A(n41403), .B(w_pixel_count[6]), 
         .C(w_pixel_count[7]), .D(n41449), .Z(n41371)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam vr_seg_line2_I_0_3_lut_rep_284_4_lut.init = 16'h8000;
    LUT4 green_leds_fixed_11__bdd_4_lut_38456 (.A(green_leds_fixed[11]), .B(green_leds_fixed[9]), 
         .C(green_leds_fixed[8]), .D(green_leds_fixed[10]), .Z(seg7_2_6__N_3439[6])) /* synthesis lut_function=(A (B+(C+!(D)))+!A !(B (C (D))+!B !(D))) */ ;
    defparam green_leds_fixed_11__bdd_4_lut_38456.init = 16'hbdee;
    LUT4 green_leds_fixed_7__bdd_4_lut (.A(green_leds_fixed[7]), .B(green_leds_fixed[5]), 
         .C(green_leds_fixed[4]), .D(green_leds_fixed[6]), .Z(seg7_1_6__N_3432[6])) /* synthesis lut_function=(A (B+(C+!(D)))+!A !(B (C (D))+!B !(D))) */ ;
    defparam green_leds_fixed_7__bdd_4_lut.init = 16'hbdee;
    FD1S3AX seg7_2_i1 (.D(seg7_2_6__N_3439[1]), .CK(w_clk_video), .Q(seg7_2[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_2_i1.GSR = "DISABLED";
    LUT4 mux_113_i1_3_lut (.A(seg7_1[0]), .B(seg7_0[0]), .C(h_seg_line0), 
         .Z(n749[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(170[3] 182[12])
    defparam mux_113_i1_3_lut.init = 16'hcaca;
    LUT4 i42_4_lut_adj_520 (.A(n41449), .B(seg7_2[0]), .C(h_seg_line2), 
         .D(n24_adj_3978), .Z(n37473)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(173[3] 182[12])
    defparam i42_4_lut_adj_520.init = 16'hcac0;
    LUT4 mux_134_i1_3_lut (.A(n1168[0]), .B(seg7_0[5]), .C(vl_seg_line0), 
         .Z(n1172[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(210[3] 222[12])
    defparam mux_134_i1_3_lut.init = 16'hcaca;
    LUT4 mux_132_i1_3_lut (.A(n565), .B(seg7_3[5]), .C(vl_seg_line3), 
         .Z(n1164[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(216[3] 222[12])
    defparam mux_132_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut (.A(n10), .B(w_line_count[4]), .C(w_line_count[6]), 
         .D(w_line_count[5]), .Z(n38805)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_4_lut.init = 16'h0020;
    LUT4 mux_176_i1_3_lut (.A(n1840[0]), .B(seg7_0[4]), .C(vl_seg_line0), 
         .Z(n1844[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(273[3] 285[12])
    defparam mux_176_i1_3_lut.init = 16'hcaca;
    LUT4 mux_174_i1_3_lut (.A(n565), .B(seg7_3[4]), .C(vl_seg_line3), 
         .Z(n1836[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(279[3] 285[12])
    defparam mux_174_i1_3_lut.init = 16'hcaca;
    LUT4 mux_197_i1_3_lut (.A(seg7_1[3]), .B(seg7_0[3]), .C(h_seg_line0), 
         .Z(n2093[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(296[3] 308[12])
    defparam mux_197_i1_3_lut.init = 16'hcaca;
    LUT4 i42_4_lut_adj_521 (.A(n41449), .B(seg7_2[3]), .C(h_seg_line2), 
         .D(n24_adj_3979), .Z(n37487)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(299[3] 308[12])
    defparam i42_4_lut_adj_521.init = 16'hcac0;
    LUT4 i1_4_lut_adj_522 (.A(n41420), .B(n25681), .C(n32490), .D(w_line_count[7]), 
         .Z(n534)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_522.init = 16'h0400;
    LUT4 green_leds_fixed_9__bdd_4_lut (.A(green_leds_fixed[9]), .B(green_leds_fixed[8]), 
         .C(green_leds_fixed[11]), .D(green_leds_fixed[10]), .Z(seg7_2_6__N_3439[5])) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A !(B (C (D)+!C !(D)))) */ ;
    defparam green_leds_fixed_9__bdd_4_lut.init = 16'hb7f1;
    LUT4 i1_4_lut_adj_523 (.A(w_line_count[3]), .B(n24402), .C(w_line_count[4]), 
         .D(n6_adj_3980), .Z(n25681)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;
    defparam i1_4_lut_adj_523.init = 16'hfcec;
    LUT4 i29909_4_lut (.A(n41511), .B(n24402), .C(w_line_count[1]), .D(w_line_count[4]), 
         .Z(n32490)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i29909_4_lut.init = 16'heccc;
    LUT4 i1_4_lut_adj_524 (.A(n41420), .B(n25680), .C(n32561), .D(w_line_count[7]), 
         .Z(n759)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_524.init = 16'h0400;
    LUT4 i1_4_lut_adj_525 (.A(w_line_count[3]), .B(n24402), .C(n6_adj_3980), 
         .D(w_line_count[4]), .Z(n25680)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_525.init = 16'heccc;
    LUT4 i21781_2_lut (.A(w_line_count[5]), .B(w_line_count[6]), .Z(n24402)) /* synthesis lut_function=(A+(B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(162[29:48])
    defparam i21781_2_lut.init = 16'heeee;
    LUT4 mux_197_i2_3_lut (.A(seg7_1[3]), .B(seg7_0[3]), .C(h_seg_line0), 
         .Z(n2093[1])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(296[3] 308[12])
    defparam mux_197_i2_3_lut.init = 16'h3535;
    LUT4 mux_180_i2_4_lut_4_lut (.A(n41383), .B(vr_seg_line3), .C(seg7_3[2]), 
         .D(n1848[1]), .Z(n1860[1])) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(201[3] 222[12])
    defparam mux_180_i2_4_lut_4_lut.init = 16'h1d0c;
    LUT4 mux_196_i2_4_lut (.A(n41369), .B(seg7_2[3]), .C(h_seg_line2), 
         .D(seg7_3[3]), .Z(n2089[1])) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(299[3] 308[12])
    defparam mux_196_i2_4_lut.init = 16'h303a;
    LUT4 mux_138_i2_4_lut_4_lut (.A(n41383), .B(vr_seg_line3), .C(seg7_3[1]), 
         .D(n1176[1]), .Z(n1188[1])) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C)+!B !(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(201[3] 222[12])
    defparam mux_138_i2_4_lut_4_lut.init = 16'h1d0c;
    LUT4 i33_4_lut_adj_526 (.A(green_leds_fixed[3]), .B(green_leds_fixed[1]), 
         .C(green_leds_fixed[0]), .D(green_leds_fixed[2]), .Z(seg7_0_6__N_3425[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D)))+!A (B (C (D))+!B !(C (D)+!C !(D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(106[2] 123[9])
    defparam i33_4_lut_adj_526.init = 16'h3ee7;
    LUT4 i38080_2_lut_2_lut_4_lut (.A(n41404), .B(n38829), .C(n38805), 
         .D(n41389), .Z(n39595)) /* synthesis lut_function=(!(A (D)+!A !(B+(C+!(D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(155[2] 311[11])
    defparam i38080_2_lut_2_lut_4_lut.init = 16'h54ff;
    LUT4 i38074_2_lut_4_lut (.A(n41404), .B(n38829), .C(n38805), .D(n534), 
         .Z(n39599)) /* synthesis lut_function=(A (D)+!A (B+(C+(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(155[2] 311[11])
    defparam i38074_2_lut_4_lut.init = 16'hff54;
    LUT4 i36858_2_lut_rep_302 (.A(n534), .B(n759), .Z(n41389)) /* synthesis lut_function=(!(A+(B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(185[2] 311[11])
    defparam i36858_2_lut_rep_302.init = 16'h1111;
    LUT4 green_leds_fixed_15__bdd_4_lut_38458 (.A(green_leds_fixed[15]), .B(green_leds_fixed[13]), 
         .C(green_leds_fixed[12]), .D(green_leds_fixed[14]), .Z(seg7_3_6__N_3446[6])) /* synthesis lut_function=(A (B+(C+!(D)))+!A !(B (C (D))+!B !(D))) */ ;
    defparam green_leds_fixed_15__bdd_4_lut_38458.init = 16'hbdee;
    PFUMX mux_177_i1 (.BLUT(n1836[0]), .ALUT(n1844[0]), .C0(n39292), .Z(n1848[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;
    LUT4 i36863_2_lut_3_lut_4_lut (.A(n534), .B(n759), .C(n38829), .D(n41404), 
         .Z(n39417)) /* synthesis lut_function=(!(A+(B+!((D)+!C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(185[2] 311[11])
    defparam i36863_2_lut_3_lut_4_lut.init = 16'h1101;
    PFUMX mux_135_i1 (.BLUT(n1164[0]), .ALUT(n1172[0]), .C0(n39292), .Z(n1176[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;
    PFUMX mux_114_i1 (.BLUT(n37473), .ALUT(n749[0]), .C0(n41358), .Z(n753[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;
    LUT4 i1_4_lut_adj_527 (.A(n41487), .B(n39164), .C(n16), .D(w_pixel_count[8]), 
         .Z(vr_seg_line1)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_527.init = 16'h1000;
    LUT4 green_leds_fixed_5__bdd_4_lut_38462 (.A(green_leds_fixed[5]), .B(green_leds_fixed[4]), 
         .C(green_leds_fixed[7]), .D(green_leds_fixed[6]), .Z(seg7_1_6__N_3432[5])) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A !(B (C (D)+!C !(D)))) */ ;
    defparam green_leds_fixed_5__bdd_4_lut_38462.init = 16'hb7f1;
    LUT4 i3_1_lut (.A(w_pixel_count[6]), .Z(led_idx[1])) /* synthesis lut_function=(!(A)) */ ;
    defparam i3_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_rep_411 (.A(w_line_count[5]), .B(w_line_count[4]), .Z(n41498)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_411.init = 16'h8888;
    LUT4 i1_4_lut_4_lut_adj_528 (.A(w_line_count[5]), .B(w_line_count[4]), 
         .C(n10), .D(w_line_count[6]), .Z(n38829)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i1_4_lut_4_lut_adj_528.init = 16'h2000;
    LUT4 i36617_2_lut (.A(w_pixel_count[7]), .B(w_pixel_count[6]), .Z(n39164)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i36617_2_lut.init = 16'heeee;
    LUT4 i29977_3_lut_4_lut (.A(w_line_count[5]), .B(w_line_count[4]), .C(w_line_count[6]), 
         .D(n41521), .Z(n32561)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;
    defparam i29977_3_lut_4_lut.init = 16'hf8f0;
    LUT4 i38069_4_lut (.A(n41420), .B(n14), .C(n32519), .D(w_line_count[7]), 
         .Z(n1431)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(248[6:48])
    defparam i38069_4_lut.init = 16'hfbff;
    LUT4 i20226_4_lut (.A(n41498), .B(w_line_count[6]), .C(n41447), .D(w_line_count[3]), 
         .Z(n14)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i20226_4_lut.init = 16'heccc;
    LUT4 mux_155_i1_3_lut (.A(n1417[0]), .B(seg7_1[6]), .C(h_seg_line1), 
         .Z(n1421[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(233[3] 245[12])
    defparam mux_155_i1_3_lut.init = 16'hcaca;
    LUT4 mux_154_i1_4_lut (.A(seg7_3[6]), .B(seg7_2[6]), .C(h_seg_line2), 
         .D(n41369), .Z(n1417[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(236[3] 245[12])
    defparam mux_154_i1_4_lut.init = 16'hcac0;
    LUT4 green_leds_fixed_3__bdd_4_lut (.A(green_leds_fixed[3]), .B(green_leds_fixed[1]), 
         .C(green_leds_fixed[0]), .D(green_leds_fixed[2]), .Z(seg7_0_6__N_3425[6])) /* synthesis lut_function=(A (B+(C+!(D)))+!A !(B (C (D))+!B !(D))) */ ;
    defparam green_leds_fixed_3__bdd_4_lut.init = 16'hbdee;
    LUT4 green_leds_fixed_1__bdd_4_lut (.A(green_leds_fixed[1]), .B(green_leds_fixed[0]), 
         .C(green_leds_fixed[3]), .D(green_leds_fixed[2]), .Z(seg7_0_6__N_3425[5])) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A !(B (C (D)+!C !(D)))) */ ;
    defparam green_leds_fixed_1__bdd_4_lut.init = 16'hb7f1;
    PFUMX mux_135_i2 (.BLUT(n1168[1]), .ALUT(n1172[1]), .C0(n39524), .Z(n1176[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;
    LUT4 i27062_4_lut (.A(n31868), .B(w_pixel_count[6]), .C(n29670), .D(w_pixel_count[7]), 
         .Z(n29675)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A (B (D)+!B !(C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(27[12:25])
    defparam i27062_4_lut.init = 16'h10fc;
    LUT4 i4_4_lut (.A(n39164), .B(n38917), .C(w_pixel_count[8]), .D(n41487), 
         .Z(h_seg_line1)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i4_4_lut.init = 16'h0040;
    LUT4 i1_4_lut_adj_529 (.A(n41420), .B(n14_adj_3981), .C(n32447), .D(w_line_count[7]), 
         .Z(n1206)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_529.init = 16'h0400;
    LUT4 i20274_3_lut (.A(n41415), .B(w_line_count[6]), .C(w_line_count[5]), 
         .Z(n14_adj_3981)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i20274_3_lut.init = 16'hecec;
    LUT4 i29873_4_lut (.A(w_line_count[2]), .B(w_line_count[6]), .C(n41520), 
         .D(w_line_count[5]), .Z(n32447)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i29873_4_lut.init = 16'heccc;
    LUT4 i20286_2_lut_rep_316_3_lut_4_lut (.A(n41518), .B(w_pixel_count[2]), 
         .C(w_pixel_count[5]), .D(n41489), .Z(n41403)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i20286_2_lut_rep_316_3_lut_4_lut.init = 16'he000;
    PFUMX mux_177_i2 (.BLUT(n1840[1]), .ALUT(n1844[1]), .C0(n39524), .Z(n1848[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;
    LUT4 mux_8_Mux_2_i15_4_lut (.A(green_leds_fixed[2]), .B(green_leds_fixed[0]), 
         .C(green_leds_fixed[3]), .D(green_leds_fixed[1]), .Z(seg7_0_6__N_3425[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A !(B+(C+!(D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(106[2] 123[9])
    defparam mux_8_Mux_2_i15_4_lut.init = 16'h5edf;
    PFUMX mux_182_i2 (.BLUT(n1864[1]), .ALUT(n1432[1]), .C0(vr_seg_line0), 
          .Z(n1868[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;
    LUT4 green_leds_fixed_5__bdd_4_lut (.A(green_leds_fixed[5]), .B(green_leds_fixed[7]), 
         .C(green_leds_fixed[6]), .D(green_leds_fixed[4]), .Z(seg7_1_6__N_3432[1])) /* synthesis lut_function=(!(A (B (C+(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C (D))))) */ ;
    defparam green_leds_fixed_5__bdd_4_lut.init = 16'h671f;
    LUT4 green_leds_fixed_11__bdd_4_lut (.A(green_leds_fixed[11]), .B(green_leds_fixed[9]), 
         .C(green_leds_fixed[8]), .D(green_leds_fixed[10]), .Z(seg7_2_6__N_3439[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D)))+!A (B (C (D))+!B !(C (D)+!C !(D))))) */ ;
    defparam green_leds_fixed_11__bdd_4_lut.init = 16'h3ee7;
    LUT4 i23384_3_lut (.A(n1431), .B(n759), .C(n1206), .Z(n26024)) /* synthesis lut_function=(A (B)+!A (B+!(C))) */ ;
    defparam i23384_3_lut.init = 16'hcdcd;
    LUT4 i2_4_lut (.A(n41371), .B(n41487), .C(n44), .D(n4_adj_3976), 
         .Z(n6)) /* synthesis lut_function=(A+!(B+!(C+(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(252[3] 285[12])
    defparam i2_4_lut.init = 16'hbbba;
    FD1S3IX color_fixed_i2 (.D(color_2__N_3467[2]), .CK(w_clk_video), .CD(n41378), 
            .Q(color_fixed[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(315[8] 316[21])
    defparam color_fixed_i2.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_530 (.A(w_pixel_count[8]), .B(n39164), .C(n4_adj_3977), 
         .D(n16), .Z(n44)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(252[3] 285[12])
    defparam i1_4_lut_adj_530.init = 16'ha2a0;
    LUT4 green_leds_fixed_15__bdd_4_lut (.A(green_leds_fixed[15]), .B(green_leds_fixed[13]), 
         .C(green_leds_fixed[12]), .D(green_leds_fixed[14]), .Z(seg7_3_6__N_3446[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D)))+!A (B (C (D))+!B !(C (D)+!C !(D))))) */ ;
    defparam green_leds_fixed_15__bdd_4_lut.init = 16'h3ee7;
    LUT4 green_leds_fixed_13__bdd_4_lut (.A(green_leds_fixed[13]), .B(green_leds_fixed[15]), 
         .C(green_leds_fixed[14]), .D(green_leds_fixed[12]), .Z(seg7_3_6__N_3446[1])) /* synthesis lut_function=(!(A (B (C+(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C (D))))) */ ;
    defparam green_leds_fixed_13__bdd_4_lut.init = 16'h671f;
    LUT4 i1_4_lut_adj_531 (.A(w_pixel_count[6]), .B(n41368), .C(w_pixel_count[8]), 
         .D(n4_adj_3982), .Z(n4_adj_3976)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_4_lut_adj_531.init = 16'h0040;
    LUT4 i1_2_lut_adj_532 (.A(w_pixel_count[5]), .B(w_pixel_count[7]), .Z(n4_adj_3982)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_532.init = 16'heeee;
    LUT4 i23387_4_lut (.A(n26020), .B(n534), .C(n26024), .D(n1206), 
         .Z(n26027)) /* synthesis lut_function=(A (B+!(C))+!A (B+!(C+!(D)))) */ ;
    defparam i23387_4_lut.init = 16'hcfce;
    LUT4 i23380_2_lut (.A(n1878), .B(n1431), .Z(n26020)) /* synthesis lut_function=(A (B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(248[2] 311[11])
    defparam i23380_2_lut.init = 16'h8888;
    FD1S3AX color_fixed_i1 (.D(color[1]), .CK(w_clk_video), .Q(color_fixed[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(315[8] 316[21])
    defparam color_fixed_i1.GSR = "DISABLED";
    LUT4 i1_4_lut_adj_533 (.A(n41420), .B(n12), .C(n32466), .D(n41522), 
         .Z(n1878)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_4_lut_adj_533.init = 16'h0400;
    LUT4 i1_4_lut_4_lut_adj_534 (.A(n41386), .B(w_pixel_count[7]), .C(w_pixel_count[8]), 
         .D(n41487), .Z(vr_seg_line0)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_4_lut_4_lut_adj_534.init = 16'h0020;
    LUT4 green_leds_fixed_0__bdd_4_lut (.A(green_leds_fixed[0]), .B(green_leds_fixed[3]), 
         .C(green_leds_fixed[2]), .D(green_leds_fixed[1]), .Z(seg7_0_6__N_3425[4])) /* synthesis lut_function=(A (B (C+(D)))+!A (B+((D)+!C))) */ ;
    defparam green_leds_fixed_0__bdd_4_lut.init = 16'hddc5;
    FD1S3AX seg7_3_i6 (.D(seg7_3_6__N_3446[6]), .CK(w_clk_video), .Q(seg7_3[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_3_i6.GSR = "DISABLED";
    FD1S3AX seg7_3_i5 (.D(seg7_3_6__N_3446[5]), .CK(w_clk_video), .Q(seg7_3[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_3_i5.GSR = "DISABLED";
    FD1S3AX seg7_3_i4 (.D(seg7_3_6__N_3446[4]), .CK(w_clk_video), .Q(seg7_3[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_3_i4.GSR = "DISABLED";
    LUT4 i37833_2_lut_rep_273_4_lut (.A(n41449), .B(n41386), .C(w_pixel_count[7]), 
         .D(vr_seg_line1), .Z(n41360)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(99[42:89])
    defparam i37833_2_lut_rep_273_4_lut.init = 16'hff80;
    FD1S3AX seg7_3_i3 (.D(seg7_3_6__N_3446[3]), .CK(w_clk_video), .Q(seg7_3[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_3_i3.GSR = "DISABLED";
    LUT4 red_leds_fixed_15__I_171_2_lut (.A(r_vsync_), .B(vsync_c), .Z(red_leds_fixed_15__N_3476)) /* synthesis lut_function=(!(A+!(B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(65[6:37])
    defparam red_leds_fixed_15__I_171_2_lut.init = 16'h4444;
    FD1S3AX seg7_3_i2 (.D(seg7_3_6__N_3446[2]), .CK(w_clk_video), .Q(seg7_3[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_3_i2.GSR = "DISABLED";
    LUT4 mux_140_i2_3_lut (.A(n1192[1]), .B(seg7_0[1]), .C(vr_seg_line0), 
         .Z(n1196[1])) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(192[3] 222[12])
    defparam mux_140_i2_3_lut.init = 16'h3a3a;
    LUT4 mux_140_i1_3_lut (.A(n1192[0]), .B(seg7_0[1]), .C(vr_seg_line0), 
         .Z(n1196[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(192[3] 222[12])
    defparam mux_140_i1_3_lut.init = 16'hcaca;
    LUT4 mux_138_i1_4_lut (.A(n1176[0]), .B(seg7_3[1]), .C(vr_seg_line3), 
         .D(n41383), .Z(n1188[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(198[3] 222[12])
    defparam mux_138_i1_4_lut.init = 16'hcfca;
    LUT4 mux_202_i1_3_lut (.A(n753[0]), .B(color_2__N_3470[0]), .C(n41388), 
         .Z(n2113[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(225[2] 311[11])
    defparam mux_202_i1_3_lut.init = 16'hcaca;
    FD1S3AX seg7_3_i1 (.D(seg7_3_6__N_3446[1]), .CK(w_clk_video), .Q(seg7_3[1])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_3_i1.GSR = "DISABLED";
    LUT4 mux_181_i1_3_lut (.A(seg7_2[2]), .B(seg7_1[2]), .C(vr_seg_line1), 
         .Z(n1864[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(258[3] 285[12])
    defparam mux_181_i1_3_lut.init = 16'hcaca;
    LUT4 mux_180_i1_4_lut (.A(n1848[0]), .B(seg7_3[2]), .C(vr_seg_line3), 
         .D(n41383), .Z(n1860[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(261[3] 285[12])
    defparam mux_180_i1_4_lut.init = 16'hcfca;
    FD1S3AX seg7_2_i6 (.D(seg7_2_6__N_3439[6]), .CK(w_clk_video), .Q(seg7_2[6])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_2_i6.GSR = "DISABLED";
    LUT4 i20170_2_lut_3_lut_4_lut (.A(n41418), .B(w_pixel_count[5]), .C(w_pixel_count[7]), 
         .D(w_pixel_count[6]), .Z(n16_adj_3983)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i20170_2_lut_3_lut_4_lut.init = 16'hfef0;
    FD1S3AX seg7_2_i5 (.D(seg7_2_6__N_3439[5]), .CK(w_clk_video), .Q(seg7_2[5])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_2_i5.GSR = "DISABLED";
    FD1S3AX seg7_2_i4 (.D(seg7_2_6__N_3439[4]), .CK(w_clk_video), .Q(seg7_2[4])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_2_i4.GSR = "DISABLED";
    FD1S3AX seg7_2_i3 (.D(seg7_2_6__N_3439[3]), .CK(w_clk_video), .Q(seg7_2[3])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_2_i3.GSR = "DISABLED";
    FD1S3AX seg7_2_i2 (.D(seg7_2_6__N_3439[2]), .CK(w_clk_video), .Q(seg7_2[2])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(134[8] 142[4])
    defparam seg7_2_i2.GSR = "DISABLED";
    LUT4 i20216_2_lut_rep_281_3_lut_4_lut (.A(n41418), .B(w_pixel_count[5]), 
         .C(w_pixel_count[7]), .D(w_pixel_count[6]), .Z(n41368)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i20216_2_lut_rep_281_3_lut_4_lut.init = 16'hfffe;
    LUT4 i20233_3_lut_4_lut (.A(n41418), .B(w_pixel_count[5]), .C(w_pixel_count[6]), 
         .D(w_pixel_count[7]), .Z(n16)) /* synthesis lut_function=(A (B+(C+(D)))+!A (C+(D))) */ ;
    defparam i20233_3_lut_4_lut.init = 16'hfff8;
    LUT4 w_pixel_count_6__bdd_3_lut_rep_296_4_lut (.A(n41418), .B(w_pixel_count[5]), 
         .C(n41449), .D(w_pixel_count[7]), .Z(n41383)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam w_pixel_count_6__bdd_3_lut_rep_296_4_lut.init = 16'h0080;
    LUT4 i2_3_lut_4_lut_adj_535 (.A(n41418), .B(w_pixel_count[5]), .C(w_pixel_count[6]), 
         .D(n41416), .Z(vr_seg_line3)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i2_3_lut_4_lut_adj_535.init = 16'h0800;
    LUT4 i36638_3_lut_rep_301_4_lut (.A(w_line_count[7]), .B(n41420), .C(n38805), 
         .D(n38829), .Z(n41388)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(155[25:41])
    defparam i36638_3_lut_rep_301_4_lut.init = 16'h1110;
    LUT4 i38076_2_lut_3_lut (.A(color_fixed[0]), .B(color_fixed[1]), .C(color_fixed[2]), 
         .Z(r_c_0)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(314[10:21])
    defparam i38076_2_lut_3_lut.init = 16'hf9f9;
    LUT4 color_fixed_2__bdd_3_lut (.A(color_fixed[2]), .B(color_fixed[0]), 
         .C(color_fixed[1]), .Z(b_c_0)) /* synthesis lut_function=(A (B (C))+!A !(B+(C))) */ ;
    defparam color_fixed_2__bdd_3_lut.init = 16'h8181;
    LUT4 green_leds_fixed_4__bdd_4_lut_38241 (.A(green_leds_fixed[4]), .B(green_leds_fixed[7]), 
         .C(green_leds_fixed[5]), .D(green_leds_fixed[6]), .Z(seg7_1_6__N_3432[0])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+(D)))+!A (B+(C+!(D)))) */ ;
    defparam green_leds_fixed_4__bdd_4_lut_38241.init = 16'hf67d;
    LUT4 green_leds_fixed_9__bdd_4_lut_38198 (.A(green_leds_fixed[9]), .B(green_leds_fixed[11]), 
         .C(green_leds_fixed[10]), .D(green_leds_fixed[8]), .Z(seg7_2_6__N_3439[1])) /* synthesis lut_function=(!(A (B (C+(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C (D))))) */ ;
    defparam green_leds_fixed_9__bdd_4_lut_38198.init = 16'h671f;
    LUT4 mux_182_i1_3_lut (.A(n1864[0]), .B(seg7_0[2]), .C(vr_seg_line0), 
         .Z(n1868[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(255[3] 285[12])
    defparam mux_182_i1_3_lut.init = 16'hcaca;
    LUT4 mux_156_i1_3_lut (.A(n1421[0]), .B(seg7_0[6]), .C(h_seg_line0), 
         .Z(n1425[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(230[3] 245[12])
    defparam mux_156_i1_3_lut.init = 16'hcaca;
    LUT4 mux_139_i1_3_lut (.A(seg7_2[1]), .B(seg7_1[1]), .C(vr_seg_line1), 
         .Z(n1192[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(195[3] 222[12])
    defparam mux_139_i1_3_lut.init = 16'hcaca;
    LUT4 mux_139_i2_3_lut (.A(seg7_2[1]), .B(seg7_1[1]), .C(vr_seg_line1), 
         .Z(n1192[1])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(195[3] 222[12])
    defparam mux_139_i2_3_lut.init = 16'h3535;
    LUT4 mux_113_i2_3_lut (.A(seg7_1[0]), .B(seg7_0[0]), .C(h_seg_line0), 
         .Z(n749[1])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(170[3] 182[12])
    defparam mux_113_i2_3_lut.init = 16'h3535;
    LUT4 mux_112_i2_4_lut (.A(seg7_3[0]), .B(seg7_2[0]), .C(h_seg_line2), 
         .D(n41369), .Z(n745[1])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(173[3] 182[12])
    defparam mux_112_i2_4_lut.init = 16'h3530;
    LUT4 i4_4_lut_adj_536 (.A(h_seg_line2), .B(h_seg_line0), .C(h_seg_line1), 
         .D(n41617), .Z(n36826)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i4_4_lut_adj_536.init = 16'hfffe;
    LUT4 i20160_2_lut_rep_314_3_lut_4_lut (.A(n41518), .B(w_pixel_count[2]), 
         .C(w_pixel_count[5]), .D(n41489), .Z(n41401)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (C))) */ ;
    defparam i20160_2_lut_rep_314_3_lut_4_lut.init = 16'hfef0;
    LUT4 green_leds_fixed_8__bdd_4_lut (.A(green_leds_fixed[8]), .B(green_leds_fixed[11]), 
         .C(green_leds_fixed[9]), .D(green_leds_fixed[10]), .Z(seg7_2_6__N_3439[0])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+(D)))+!A (B+(C+!(D)))) */ ;
    defparam green_leds_fixed_8__bdd_4_lut.init = 16'hf67d;
    L6MUX21 i37241 (.D0(n39793), .D1(n39794), .SD(w_pixel_count[8]), .Z(color_2__N_3479[0]));
    LUT4 i1_2_lut_rep_282_3_lut_4_lut (.A(w_pixel_count[8]), .B(n41487), 
         .C(n29675), .D(w_pixel_count[7]), .Z(n41369)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(173[3] 182[12])
    defparam i1_2_lut_rep_282_3_lut_4_lut.init = 16'h1000;
    LUT4 h_seg_line0_I_0_4_lut_4_lut_4_lut (.A(w_pixel_count[8]), .B(n41487), 
         .C(n36829), .D(n213), .Z(h_seg_line0)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C)+!B !(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(173[3] 182[12])
    defparam h_seg_line0_I_0_4_lut_4_lut_4_lut.init = 16'h1f0c;
    LUT4 green_leds_fixed_0__bdd_4_lut_38451 (.A(green_leds_fixed[0]), .B(green_leds_fixed[3]), 
         .C(green_leds_fixed[1]), .D(green_leds_fixed[2]), .Z(seg7_0_6__N_3425[0])) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C+(D)))+!A (B+(C+!(D)))) */ ;
    defparam green_leds_fixed_0__bdd_4_lut_38451.init = 16'hf67d;
    LUT4 i37228_3_lut_3_lut (.A(w_pixel_count[5]), .B(green_leds_fixed[11]), 
         .C(green_leds_fixed[10]), .Z(n39782)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(78[37:70])
    defparam i37228_3_lut_3_lut.init = 16'he4e4;
    LUT4 i37227_3_lut_3_lut (.A(w_pixel_count[5]), .B(green_leds_fixed[9]), 
         .C(green_leds_fixed[8]), .Z(n39781)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(78[37:70])
    defparam i37227_3_lut_3_lut.init = 16'he4e4;
    LUT4 green_leds_fixed_1__bdd_4_lut_38429 (.A(green_leds_fixed[1]), .B(green_leds_fixed[3]), 
         .C(green_leds_fixed[2]), .D(green_leds_fixed[0]), .Z(seg7_0_6__N_3425[1])) /* synthesis lut_function=(!(A (B (C+(D))+!B !((D)+!C))+!A !(B ((D)+!C)+!B !(C (D))))) */ ;
    defparam green_leds_fixed_1__bdd_4_lut_38429.init = 16'h671f;
    FD1P3AX green_leds_fixed_i0_i0 (.D(\counter[0] ), .SP(red_leds_fixed_15__N_3476), 
            .CK(w_clk_video), .Q(green_leds_fixed[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=47, LSE_RLINE=58 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(59[8] 71[4])
    defparam green_leds_fixed_i0_i0.GSR = "DISABLED";
    LUT4 i37231_3_lut_3_lut (.A(w_pixel_count[5]), .B(green_leds_fixed[1]), 
         .C(green_leds_fixed[0]), .Z(n39785)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(78[37:70])
    defparam i37231_3_lut_3_lut.init = 16'he4e4;
    LUT4 i37230_3_lut_3_lut (.A(w_pixel_count[5]), .B(green_leds_fixed[15]), 
         .C(green_leds_fixed[14]), .Z(n39784)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(78[37:70])
    defparam i37230_3_lut_3_lut.init = 16'he4e4;
    LUT4 i37233_3_lut_3_lut (.A(w_pixel_count[5]), .B(green_leds_fixed[5]), 
         .C(green_leds_fixed[4]), .Z(n39787)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(78[37:70])
    defparam i37233_3_lut_3_lut.init = 16'he4e4;
    LUT4 i37229_3_lut_3_lut (.A(w_pixel_count[5]), .B(green_leds_fixed[13]), 
         .C(green_leds_fixed[12]), .Z(n39783)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(78[37:70])
    defparam i37229_3_lut_3_lut.init = 16'he4e4;
    LUT4 i1_2_lut_rep_400 (.A(w_pixel_count[10]), .B(w_pixel_count[9]), 
         .Z(n41487)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_400.init = 16'heeee;
    LUT4 i1_2_lut_rep_329_3_lut_4_lut (.A(w_pixel_count[10]), .B(w_pixel_count[9]), 
         .C(w_pixel_count[7]), .D(w_pixel_count[8]), .Z(n41416)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i1_2_lut_rep_329_3_lut_4_lut.init = 16'h0010;
    LUT4 i37879_2_lut_rep_362_3_lut (.A(w_pixel_count[10]), .B(w_pixel_count[9]), 
         .C(w_pixel_count[8]), .Z(n41449)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i37879_2_lut_rep_362_3_lut.init = 16'h0101;
    LUT4 mux_202_i2_3_lut_4_lut (.A(n41404), .B(n38805), .C(color_2__N_3470[1]), 
         .D(n745[1]), .Z(n2113[1])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_202_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 i38088_2_lut_3_lut_4_lut (.A(w_pixel_count[10]), .B(w_pixel_count[9]), 
         .C(vl_seg_line0), .D(n4_adj_3976), .Z(n39524)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i38088_2_lut_3_lut_4_lut.init = 16'hf1f0;
    LUT4 b_c_bdd_2_lut_38197_3_lut_4_lut (.A(w_pixel_count[10]), .B(w_pixel_count[9]), 
         .C(n40635), .D(w_pixel_count[8]), .Z(n40636)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam b_c_bdd_2_lut_38197_3_lut_4_lut.init = 16'h0010;
    LUT4 mux_114_i2_3_lut_4_lut (.A(n41404), .B(n38829), .C(color_2__N_3470[0]), 
         .D(n749[1]), .Z(n753[1])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam mux_114_i2_3_lut_4_lut.init = 16'hfb40;
    LUT4 i20168_1_lut_rep_389 (.A(w_pixel_count[7]), .Z(n41476)) /* synthesis lut_function=(!(A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(91[42:65])
    defparam i20168_1_lut_rep_389.init = 16'h5555;
    LUT4 i1_4_lut_4_lut_adj_537 (.A(w_pixel_count[7]), .B(n4_adj_3984), 
         .C(n4_adj_3977), .D(n41449), .Z(n565)) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(91[42:65])
    defparam i1_4_lut_4_lut_adj_537.init = 16'hf400;
    LUT4 i37830_2_lut_3_lut_4_lut_4_lut (.A(n41404), .B(n38829), .C(n534), 
         .D(n38805), .Z(n39428)) /* synthesis lut_function=(A (C)+!A (B+(C+(D)))) */ ;
    defparam i37830_2_lut_3_lut_4_lut_4_lut.init = 16'hf5f4;
    LUT4 color_2__I_173_i3_3_lut_4_lut (.A(n41404), .B(n38829), .C(color_2__N_3470[1]), 
         .D(color_2__N_3482[2]), .Z(color_2__N_3467[2])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;
    defparam color_2__I_173_i3_3_lut_4_lut.init = 16'hfb40;
    LUT4 vr_seg_line2_N_3586_bdd_4_lut_38203 (.A(w_pixel_count[7]), .B(n41418), 
         .C(w_pixel_count[5]), .D(w_pixel_count[6]), .Z(n40635)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A !(B))) */ ;
    defparam vr_seg_line2_N_3586_bdd_4_lut_38203.init = 16'h4ccc;
    LUT4 i1_2_lut_rep_402 (.A(w_pixel_count[4]), .B(w_pixel_count[3]), .Z(n41489)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_402.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_538 (.A(w_pixel_count[4]), .B(w_pixel_count[3]), 
         .C(w_pixel_count[5]), .Z(n31868)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_538.init = 16'h8080;
    LUT4 i43_4_lut_adj_539 (.A(n22), .B(n29675), .C(w_pixel_count[7]), 
         .D(seg7_3[3]), .Z(n24_adj_3979)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(299[3] 308[12])
    defparam i43_4_lut_adj_539.init = 16'hca0a;
    LUT4 i1_4_lut_adj_540 (.A(n41449), .B(w_pixel_count[7]), .C(n41382), 
         .D(n41517), .Z(vl_seg_line3)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_4_lut_adj_540.init = 16'h0080;
    LUT4 i1_4_lut_adj_541 (.A(n41487), .B(n202), .C(n16_adj_3983), .D(w_pixel_count[8]), 
         .Z(vl_seg_line0)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_541.init = 16'h1000;
    LUT4 i1_4_lut_adj_542 (.A(n41449), .B(w_pixel_count[7]), .C(n41381), 
         .D(n41519), .Z(vl_seg_line2)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_4_lut_adj_542.init = 16'h0080;
    LUT4 i43_4_lut_adj_543 (.A(n22), .B(n29675), .C(w_pixel_count[7]), 
         .D(seg7_3[0]), .Z(n24_adj_3978)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(173[3] 182[12])
    defparam i43_4_lut_adj_543.init = 16'hca0a;
    LUT4 i29415_2_lut_4_lut (.A(w_pixel_count[10]), .B(w_pixel_count[9]), 
         .C(w_pixel_count[4]), .D(color_2__N_3479[0]), .Z(color_2__N_3470[1])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i29415_2_lut_4_lut.init = 16'h0010;
    LUT4 i28817_2_lut_4_lut (.A(w_pixel_count[10]), .B(w_pixel_count[9]), 
         .C(w_pixel_count[4]), .D(color_2__N_3479[0]), .Z(color_2__N_3470[0])) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i28817_2_lut_4_lut.init = 16'h1000;
    PFUMX i37235 (.BLUT(n39781), .ALUT(n39782), .C0(led_idx[1]), .Z(n39789));
    PFUMX i37236 (.BLUT(n39783), .ALUT(n39784), .C0(led_idx[1]), .Z(n39790));
    PFUMX i37237 (.BLUT(n39785), .ALUT(n39786), .C0(led_idx[1]), .Z(n39791));
    LUT4 i37232_3_lut_3_lut (.A(w_pixel_count[5]), .B(green_leds_fixed[3]), 
         .C(green_leds_fixed[2]), .Z(n39786)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(78[37:70])
    defparam i37232_3_lut_3_lut.init = 16'he4e4;
    PFUMX i37238 (.BLUT(n39787), .ALUT(n39788), .C0(led_idx[1]), .Z(n39792));
    hvsync u_hvsync (.\w_pixel_count[6] (w_pixel_count[6]), .\w_pixel_count[5] (w_pixel_count[5]), 
           .n41517(n41517), .\w_pixel_count[7] (w_pixel_count[7]), .n41401(n41401), 
           .n4(n4_adj_3984), .w_line_count({Open_0, Open_1, Open_2, 
           Open_3, w_line_count[7:6], Open_4, w_line_count[4:2], Open_5, 
           Open_6}), .n41520(n41520), .n41521(n41521), .n10(n10), .n41522(n41522), 
           .n41420(n41420), .\w_line_count[1] (w_line_count[1]), .n41447(n41447), 
           .w_vsync(w_vsync), .w_hsync(w_hsync), .reset_n_N_45(reset_n_N_45), 
           .w_clk_video(w_clk_video), .\w_line_count[5] (w_line_count[5]), 
           .\w_pixel_count[10] (w_pixel_count[10]), .\w_pixel_count[8] (w_pixel_count[8]), 
           .\w_pixel_count[9] (w_pixel_count[9]), .n32565(n32565), .\w_pixel_count[3] (w_pixel_count[3]), 
           .n41519(n41519), .\w_pixel_count[4] (w_pixel_count[4]), .n4_adj_102(n4), 
           .\w_pixel_count[0] (w_pixel_count[0]), .n6(n6_adj_3980), .n38829(n38829), 
           .n41379(n41379), .n38805(n38805), .n41378(n41378), .n29675(n29675), 
           .n38917(n38917), .n31868(n31868), .n41487(n41487), .n36829(n36829), 
           .n29670(n29670), .n213(n213), .n41415(n41415), .GND_net(GND_net), 
           .\w_pixel_count[2] (w_pixel_count[2]), .n41511(n41511), .\w_pixel_count[1] (w_pixel_count[1]), 
           .n41404(n41404), .n32519(n32519), .n32466(n32466), .n41617(n41617)) /* synthesis syn_module_defined=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(38[8] 49[3])
    
endmodule
//
// Verilog Description of module hvsync
//

module hvsync (\w_pixel_count[6] , \w_pixel_count[5] , n41517, \w_pixel_count[7] , 
            n41401, n4, w_line_count, n41520, n41521, n10, n41522, 
            n41420, \w_line_count[1] , n41447, w_vsync, w_hsync, reset_n_N_45, 
            w_clk_video, \w_line_count[5] , \w_pixel_count[10] , \w_pixel_count[8] , 
            \w_pixel_count[9] , n32565, \w_pixel_count[3] , n41519, 
            \w_pixel_count[4] , n4_adj_102, \w_pixel_count[0] , n6, 
            n38829, n41379, n38805, n41378, n29675, n38917, n31868, 
            n41487, n36829, n29670, n213, n41415, GND_net, \w_pixel_count[2] , 
            n41511, \w_pixel_count[1] , n41404, n32519, n32466, n41617) /* synthesis syn_module_defined=1 */ ;
    output \w_pixel_count[6] ;
    output \w_pixel_count[5] ;
    output n41517;
    output \w_pixel_count[7] ;
    input n41401;
    output n4;
    output [11:0]w_line_count;
    output n41520;
    output n41521;
    output n10;
    output n41522;
    output n41420;
    output \w_line_count[1] ;
    output n41447;
    output w_vsync;
    output w_hsync;
    input reset_n_N_45;
    input w_clk_video;
    output \w_line_count[5] ;
    output \w_pixel_count[10] ;
    output \w_pixel_count[8] ;
    output \w_pixel_count[9] ;
    input n32565;
    output \w_pixel_count[3] ;
    input n41519;
    output \w_pixel_count[4] ;
    input n4_adj_102;
    output \w_pixel_count[0] ;
    output n6;
    input n38829;
    output n41379;
    input n38805;
    output n41378;
    input n29675;
    input n38917;
    input n31868;
    input n41487;
    output n36829;
    input n29670;
    output n213;
    output n41415;
    input GND_net;
    output \w_pixel_count[2] ;
    output n41511;
    output \w_pixel_count[1] ;
    output n41404;
    output n32519;
    output n32466;
    output n41617;
    
    wire w_hsync /* synthesis is_clock=1, SET_AS_NETWORK=\r_3__I_0/w_hsync */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(24[6:13])
    wire w_clk_video /* synthesis SET_AS_NETWORK=w_clk_video, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(21[6:17])
    
    wire n41524, n41468;
    wire [11:0]w_line_count_c;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(28[12:24])
    
    wire n41523, n41465, n39060, n38922, n11, vsync_N_3645, hsync_N_3642, 
        n39197;
    wire [11:0]n26;
    
    wire n38821, n38937, n32575;
    wire [11:0]line_count_11__N_3629;
    
    wire n38869;
    wire [10:0]n49;
    
    wire n36735;
    wire [10:0]n62;
    
    wire n41616, n41615, n36619, n36618, n36617, n36616, n36615, 
        n36614, n4_adj_3975, n36844, n36657, n36656, n36655, n36654, 
        n36653;
    
    LUT4 i1_2_lut_rep_430 (.A(\w_pixel_count[6] ), .B(\w_pixel_count[5] ), 
         .Z(n41517)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_430.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(\w_pixel_count[6] ), .B(\w_pixel_count[5] ), 
         .C(\w_pixel_count[7] ), .D(n41401), .Z(n4)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h1110;
    LUT4 i29296_2_lut_rep_433 (.A(w_line_count[3]), .B(w_line_count[4]), 
         .Z(n41520)) /* synthesis lut_function=(A (B)) */ ;
    defparam i29296_2_lut_rep_433.init = 16'h8888;
    LUT4 i1_2_lut_rep_434 (.A(w_line_count[3]), .B(w_line_count[2]), .Z(n41521)) /* synthesis lut_function=(A+(B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam i1_2_lut_rep_434.init = 16'heeee;
    LUT4 i2_3_lut_4_lut (.A(w_line_count[3]), .B(w_line_count[2]), .C(w_line_count[4]), 
         .D(n41524), .Z(n10)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam i2_3_lut_4_lut.init = 16'hfffe;
    LUT4 i20179_2_lut_rep_381_3_lut (.A(w_line_count[3]), .B(w_line_count[2]), 
         .C(w_line_count[4]), .Z(n41468)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam i20179_2_lut_rep_381_3_lut.init = 16'he0e0;
    LUT4 i1_2_lut_rep_435 (.A(w_line_count[6]), .B(w_line_count[7]), .Z(n41522)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_435.init = 16'h8888;
    LUT4 i21629_2_lut_rep_436 (.A(w_line_count_c[10]), .B(w_line_count_c[11]), 
         .Z(n41523)) /* synthesis lut_function=(A+(B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(55[68:129])
    defparam i21629_2_lut_rep_436.init = 16'heeee;
    LUT4 i1_2_lut_rep_378_3_lut (.A(w_line_count_c[10]), .B(w_line_count_c[11]), 
         .C(w_line_count_c[9]), .Z(n41465)) /* synthesis lut_function=(A+(B+(C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(55[68:129])
    defparam i1_2_lut_rep_378_3_lut.init = 16'hfefe;
    LUT4 i36517_2_lut_3_lut (.A(w_line_count_c[10]), .B(w_line_count_c[11]), 
         .C(w_line_count_c[8]), .Z(n39060)) /* synthesis lut_function=(A+(B+(C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(55[68:129])
    defparam i36517_2_lut_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_333_3_lut_4_lut (.A(w_line_count_c[10]), .B(w_line_count_c[11]), 
         .C(w_line_count_c[8]), .D(w_line_count_c[9]), .Z(n41420)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(55[68:129])
    defparam i1_2_lut_rep_333_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_437 (.A(\w_line_count[1] ), .B(w_line_count_c[0]), 
         .Z(n41524)) /* synthesis lut_function=(A+(B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(28[12:24])
    defparam i1_2_lut_rep_437.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\w_line_count[1] ), .B(w_line_count_c[0]), 
         .C(w_line_count[3]), .D(w_line_count[2]), .Z(n38922)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(28[12:24])
    defparam i1_2_lut_3_lut_4_lut.init = 16'he000;
    LUT4 i1_2_lut_rep_360_3_lut (.A(\w_line_count[1] ), .B(w_line_count_c[0]), 
         .C(w_line_count[2]), .Z(n41447)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(28[12:24])
    defparam i1_2_lut_rep_360_3_lut.init = 16'he0e0;
    LUT4 i2_4_lut (.A(n41522), .B(w_line_count_c[9]), .C(n11), .D(n39060), 
         .Z(vsync_N_3645)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_4_lut.init = 16'h0080;
    FD1S3DX vsync_27 (.D(vsync_N_3645), .CK(w_hsync), .CD(reset_n_N_45), 
            .Q(w_vsync)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=38, LSE_RLINE=49 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam vsync_27.GSR = "DISABLED";
    FD1S3DX hsync_25 (.D(hsync_N_3642), .CK(w_clk_video), .CD(reset_n_N_45), 
            .Q(w_hsync)) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=38, LSE_RLINE=49 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(38[2] 45[5])
    defparam hsync_25.GSR = "DISABLED";
    LUT4 i22_4_lut (.A(n39197), .B(n41522), .C(\w_line_count[5] ), .D(n41468), 
         .Z(n11)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;
    defparam i22_4_lut.init = 16'h3530;
    FD1S3DX line_count__i0 (.D(n26[0]), .CK(w_hsync), .CD(reset_n_N_45), 
            .Q(w_line_count_c[0])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=38, LSE_RLINE=49 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam line_count__i0.GSR = "DISABLED";
    LUT4 i3_4_lut (.A(\w_pixel_count[10] ), .B(\w_pixel_count[8] ), .C(\w_pixel_count[9] ), 
         .D(n38821), .Z(hsync_N_3642)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(39[12:129])
    defparam i3_4_lut.init = 16'h0800;
    LUT4 i1_4_lut (.A(n32565), .B(n38937), .C(\w_pixel_count[8] ), .D(\w_pixel_count[7] ), 
         .Z(n38821)) /* synthesis lut_function=(!(A (B (C (D))+!B (C+!(D)))+!A !(B+(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(39[12:129])
    defparam i1_4_lut.init = 16'h5fcc;
    LUT4 i1_4_lut_adj_507 (.A(\w_pixel_count[3] ), .B(n41519), .C(\w_pixel_count[4] ), 
         .D(n4_adj_102), .Z(n38937)) /* synthesis lut_function=(A (B (C+(D)))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(39[12:129])
    defparam i1_4_lut_adj_507.init = 16'hc8c0;
    FD1S3DX line_count__i11 (.D(n26[11]), .CK(w_hsync), .CD(reset_n_N_45), 
            .Q(w_line_count_c[11])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=38, LSE_RLINE=49 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam line_count__i11.GSR = "DISABLED";
    FD1S3DX line_count__i10 (.D(n26[10]), .CK(w_hsync), .CD(reset_n_N_45), 
            .Q(w_line_count_c[10])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=38, LSE_RLINE=49 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam line_count__i10.GSR = "DISABLED";
    FD1S3BX line_count__i9 (.D(n26[9]), .CK(w_hsync), .PD(reset_n_N_45), 
            .Q(w_line_count_c[9])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=38, LSE_RLINE=49 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam line_count__i9.GSR = "DISABLED";
    FD1S3DX line_count__i8 (.D(n26[8]), .CK(w_hsync), .CD(reset_n_N_45), 
            .Q(w_line_count_c[8])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=38, LSE_RLINE=49 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam line_count__i8.GSR = "DISABLED";
    FD1S3BX line_count__i7 (.D(n26[7]), .CK(w_hsync), .PD(reset_n_N_45), 
            .Q(w_line_count[7])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=38, LSE_RLINE=49 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam line_count__i7.GSR = "DISABLED";
    FD1S3BX line_count__i6 (.D(n26[6]), .CK(w_hsync), .PD(reset_n_N_45), 
            .Q(w_line_count[6])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=38, LSE_RLINE=49 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam line_count__i6.GSR = "DISABLED";
    FD1S3DX line_count__i5 (.D(n26[5]), .CK(w_hsync), .CD(reset_n_N_45), 
            .Q(\w_line_count[5] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=38, LSE_RLINE=49 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam line_count__i5.GSR = "DISABLED";
    FD1S3BX line_count__i4 (.D(n26[4]), .CK(w_hsync), .PD(reset_n_N_45), 
            .Q(w_line_count[4])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=38, LSE_RLINE=49 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam line_count__i4.GSR = "DISABLED";
    FD1S3DX line_count__i3 (.D(n26[3]), .CK(w_hsync), .CD(reset_n_N_45), 
            .Q(w_line_count[3])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=38, LSE_RLINE=49 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam line_count__i3.GSR = "DISABLED";
    FD1S3DX line_count__i2 (.D(n26[2]), .CK(w_hsync), .CD(reset_n_N_45), 
            .Q(w_line_count[2])) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=38, LSE_RLINE=49 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam line_count__i2.GSR = "DISABLED";
    FD1S3DX line_count__i1 (.D(n26[1]), .CK(w_hsync), .CD(reset_n_N_45), 
            .Q(\w_line_count[1] )) /* synthesis LSE_LINE_FILE_ID=4, LSE_LCOL=8, LSE_RCOL=3, LSE_LLINE=38, LSE_RLINE=49 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam line_count__i1.GSR = "DISABLED";
    LUT4 i1_2_lut (.A(n32575), .B(line_count_11__N_3629[0]), .Z(n26[0])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut.init = 16'h4444;
    LUT4 i2_4_lut_adj_508 (.A(n41522), .B(w_line_count[4]), .C(\w_line_count[5] ), 
         .D(n38922), .Z(n38869)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_508.init = 16'ha080;
    LUT4 i29409_2_lut (.A(n49[10]), .B(n36735), .Z(n62[10])) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam i29409_2_lut.init = 16'h2222;
    LUT4 i29417_2_lut (.A(n49[9]), .B(n36735), .Z(n62[9])) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam i29417_2_lut.init = 16'h2222;
    LUT4 i29423_2_lut (.A(n49[8]), .B(n36735), .Z(n62[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam i29423_2_lut.init = 16'h2222;
    LUT4 i29424_2_lut (.A(n49[7]), .B(n36735), .Z(n62[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam i29424_2_lut.init = 16'h2222;
    LUT4 i29430_2_lut (.A(n49[6]), .B(n36735), .Z(n62[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam i29430_2_lut.init = 16'h2222;
    LUT4 i29431_2_lut (.A(n49[5]), .B(n36735), .Z(n62[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam i29431_2_lut.init = 16'h2222;
    LUT4 i29434_2_lut (.A(n49[4]), .B(n36735), .Z(n62[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam i29434_2_lut.init = 16'h2222;
    LUT4 i29435_2_lut (.A(n49[3]), .B(n36735), .Z(n62[3])) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam i29435_2_lut.init = 16'h2222;
    LUT4 i29442_2_lut (.A(n49[2]), .B(n36735), .Z(n62[2])) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam i29442_2_lut.init = 16'h2222;
    LUT4 i29443_2_lut (.A(n49[1]), .B(n36735), .Z(n62[1])) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam i29443_2_lut.init = 16'h2222;
    FD1S3DX pixel_count_19667_19668__i1 (.D(n62[0]), .CK(w_clk_video), .CD(reset_n_N_45), 
            .Q(\w_pixel_count[0] )) /* synthesis syn_use_carry_chain=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam pixel_count_19667_19668__i1.GSR = "DISABLED";
    LUT4 i28867_2_lut (.A(line_count_11__N_3629[11]), .B(n32575), .Z(n26[11])) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam i28867_2_lut.init = 16'h2222;
    LUT4 i28868_2_lut (.A(line_count_11__N_3629[10]), .B(n32575), .Z(n26[10])) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam i28868_2_lut.init = 16'h2222;
    LUT4 i28952_2_lut (.A(line_count_11__N_3629[9]), .B(n32575), .Z(n26[9])) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam i28952_2_lut.init = 16'h2222;
    LUT4 i28954_2_lut (.A(line_count_11__N_3629[8]), .B(n32575), .Z(n26[8])) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam i28954_2_lut.init = 16'h2222;
    LUT4 i28955_2_lut (.A(line_count_11__N_3629[7]), .B(n32575), .Z(n26[7])) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam i28955_2_lut.init = 16'h2222;
    LUT4 i28956_2_lut (.A(line_count_11__N_3629[6]), .B(n32575), .Z(n26[6])) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam i28956_2_lut.init = 16'h2222;
    LUT4 i28957_2_lut (.A(line_count_11__N_3629[5]), .B(n32575), .Z(n26[5])) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam i28957_2_lut.init = 16'h2222;
    LUT4 i28958_2_lut (.A(line_count_11__N_3629[4]), .B(n32575), .Z(n26[4])) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam i28958_2_lut.init = 16'h2222;
    LUT4 i1_2_lut_adj_509 (.A(n32575), .B(line_count_11__N_3629[3]), .Z(n26[3])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_509.init = 16'h4444;
    LUT4 i1_2_lut_adj_510 (.A(n32575), .B(line_count_11__N_3629[2]), .Z(n26[2])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_510.init = 16'h4444;
    LUT4 i1_2_lut_adj_511 (.A(n32575), .B(line_count_11__N_3629[1]), .Z(n26[1])) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_511.init = 16'h4444;
    LUT4 i2_3_lut (.A(w_line_count[2]), .B(w_line_count_c[0]), .C(\w_line_count[1] ), 
         .Z(n6)) /* synthesis lut_function=(A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_292_3_lut_4_lut (.A(w_line_count_c[8]), .B(n41465), 
         .C(n38829), .D(w_line_count[7]), .Z(n41379)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam i1_2_lut_rep_292_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_rep_291_3_lut_4_lut (.A(w_line_count_c[8]), .B(n41465), 
         .C(n38805), .D(w_line_count[7]), .Z(n41378)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(54[2] 61[5])
    defparam i1_2_lut_rep_291_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_3_lut_4_lut_then_4_lut (.A(n29675), .B(\w_pixel_count[8] ), 
         .C(\w_pixel_count[9] ), .D(\w_pixel_count[10] ), .Z(n41616)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam i1_3_lut_4_lut_then_4_lut.init = 16'h0002;
    LUT4 i1_3_lut_4_lut_else_4_lut (.A(n38917), .B(\w_pixel_count[8] ), 
         .C(\w_pixel_count[9] ), .D(\w_pixel_count[10] ), .Z(n41615)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam i1_3_lut_4_lut_else_4_lut.init = 16'h0002;
    LUT4 i2_4_lut_adj_512 (.A(\w_pixel_count[6] ), .B(\w_pixel_count[7] ), 
         .C(n31868), .D(n41487), .Z(n36829)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;
    defparam i2_4_lut_adj_512.init = 16'hffec;
    LUT4 i1_4_lut_adj_513 (.A(\w_pixel_count[8] ), .B(\w_pixel_count[7] ), 
         .C(\w_pixel_count[6] ), .D(n29670), .Z(n213)) /* synthesis lut_function=(A (B+(C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam i1_4_lut_adj_513.init = 16'ha888;
    LUT4 i20281_3_lut_rep_328_4_lut (.A(n41524), .B(w_line_count[2]), .C(w_line_count[4]), 
         .D(w_line_count[3]), .Z(n41415)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/display.v(28[12:24])
    defparam i20281_3_lut_rep_328_4_lut.init = 16'hf080;
    CCU2D add_15_13 (.A0(w_line_count_c[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n36619), .S0(line_count_11__N_3629[11]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(58[18:35])
    defparam add_15_13.INIT0 = 16'h5aaa;
    defparam add_15_13.INIT1 = 16'h0000;
    defparam add_15_13.INJECT1_0 = "NO";
    defparam add_15_13.INJECT1_1 = "NO";
    CCU2D add_15_11 (.A0(w_line_count_c[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(w_line_count_c[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n36618), .COUT(n36619), .S0(line_count_11__N_3629[9]), 
          .S1(line_count_11__N_3629[10]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(58[18:35])
    defparam add_15_11.INIT0 = 16'h5aaa;
    defparam add_15_11.INIT1 = 16'h5aaa;
    defparam add_15_11.INJECT1_0 = "NO";
    defparam add_15_11.INJECT1_1 = "NO";
    CCU2D add_15_9 (.A0(w_line_count[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(w_line_count_c[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n36617), .COUT(n36618), .S0(line_count_11__N_3629[7]), 
          .S1(line_count_11__N_3629[8]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(58[18:35])
    defparam add_15_9.INIT0 = 16'h5aaa;
    defparam add_15_9.INIT1 = 16'h5aaa;
    defparam add_15_9.INJECT1_0 = "NO";
    defparam add_15_9.INJECT1_1 = "NO";
    CCU2D add_15_7 (.A0(\w_line_count[5] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(w_line_count[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n36616), .COUT(n36617), .S0(line_count_11__N_3629[5]), 
          .S1(line_count_11__N_3629[6]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(58[18:35])
    defparam add_15_7.INIT0 = 16'h5aaa;
    defparam add_15_7.INIT1 = 16'h5aaa;
    defparam add_15_7.INJECT1_0 = "NO";
    defparam add_15_7.INJECT1_1 = "NO";
    CCU2D add_15_5 (.A0(w_line_count[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(w_line_count[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n36615), .COUT(n36616), .S0(line_count_11__N_3629[3]), 
          .S1(line_count_11__N_3629[4]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(58[18:35])
    defparam add_15_5.INIT0 = 16'h5aaa;
    defparam add_15_5.INIT1 = 16'h5aaa;
    defparam add_15_5.INJECT1_0 = "NO";
    defparam add_15_5.INJECT1_1 = "NO";
    CCU2D add_15_3 (.A0(\w_line_count[1] ), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(w_line_count[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n36614), .COUT(n36615), .S0(line_count_11__N_3629[1]), 
          .S1(line_count_11__N_3629[2]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(58[18:35])
    defparam add_15_3.INIT0 = 16'h5aaa;
    defparam add_15_3.INIT1 = 16'h5aaa;
    defparam add_15_3.INJECT1_0 = "NO";
    defparam add_15_3.INJECT1_1 = "NO";
    FD1S3DX pixel_count_19667_19668__i11 (.D(n62[10]), .CK(w_clk_video), 
            .CD(reset_n_N_45), .Q(\w_pixel_count[10] )) /* synthesis syn_use_carry_chain=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam pixel_count_19667_19668__i11.GSR = "DISABLED";
    FD1S3DX pixel_count_19667_19668__i10 (.D(n62[9]), .CK(w_clk_video), 
            .CD(reset_n_N_45), .Q(\w_pixel_count[9] )) /* synthesis syn_use_carry_chain=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam pixel_count_19667_19668__i10.GSR = "DISABLED";
    CCU2D add_15_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(w_line_count_c[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n36614), .S1(line_count_11__N_3629[0]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(58[18:35])
    defparam add_15_1.INIT0 = 16'hF000;
    defparam add_15_1.INIT1 = 16'h5555;
    defparam add_15_1.INJECT1_0 = "NO";
    defparam add_15_1.INJECT1_1 = "NO";
    FD1S3DX pixel_count_19667_19668__i9 (.D(n62[8]), .CK(w_clk_video), .CD(reset_n_N_45), 
            .Q(\w_pixel_count[8] )) /* synthesis syn_use_carry_chain=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam pixel_count_19667_19668__i9.GSR = "DISABLED";
    FD1S3DX pixel_count_19667_19668__i8 (.D(n62[7]), .CK(w_clk_video), .CD(reset_n_N_45), 
            .Q(\w_pixel_count[7] )) /* synthesis syn_use_carry_chain=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam pixel_count_19667_19668__i8.GSR = "DISABLED";
    FD1S3DX pixel_count_19667_19668__i7 (.D(n62[6]), .CK(w_clk_video), .CD(reset_n_N_45), 
            .Q(\w_pixel_count[6] )) /* synthesis syn_use_carry_chain=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam pixel_count_19667_19668__i7.GSR = "DISABLED";
    FD1S3DX pixel_count_19667_19668__i6 (.D(n62[5]), .CK(w_clk_video), .CD(reset_n_N_45), 
            .Q(\w_pixel_count[5] )) /* synthesis syn_use_carry_chain=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam pixel_count_19667_19668__i6.GSR = "DISABLED";
    FD1S3DX pixel_count_19667_19668__i5 (.D(n62[4]), .CK(w_clk_video), .CD(reset_n_N_45), 
            .Q(\w_pixel_count[4] )) /* synthesis syn_use_carry_chain=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam pixel_count_19667_19668__i5.GSR = "DISABLED";
    FD1S3DX pixel_count_19667_19668__i4 (.D(n62[3]), .CK(w_clk_video), .CD(reset_n_N_45), 
            .Q(\w_pixel_count[3] )) /* synthesis syn_use_carry_chain=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam pixel_count_19667_19668__i4.GSR = "DISABLED";
    FD1S3DX pixel_count_19667_19668__i3 (.D(n62[2]), .CK(w_clk_video), .CD(reset_n_N_45), 
            .Q(\w_pixel_count[2] )) /* synthesis syn_use_carry_chain=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam pixel_count_19667_19668__i3.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_424 (.A(w_line_count[2]), .B(w_line_count[3]), .Z(n41511)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_424.init = 16'h8888;
    FD1S3DX pixel_count_19667_19668__i2 (.D(n62[1]), .CK(w_clk_video), .CD(reset_n_N_45), 
            .Q(\w_pixel_count[1] )) /* synthesis syn_use_carry_chain=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam pixel_count_19667_19668__i2.GSR = "DISABLED";
    LUT4 i29162_2_lut (.A(n49[0]), .B(n36735), .Z(n62[0])) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam i29162_2_lut.init = 16'h2222;
    LUT4 i2_4_lut_adj_514 (.A(\w_pixel_count[10] ), .B(\w_pixel_count[8] ), 
         .C(\w_pixel_count[9] ), .D(n4_adj_3975), .Z(n36735)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_514.init = 16'ha080;
    LUT4 i1_4_lut_adj_515 (.A(n41519), .B(\w_pixel_count[7] ), .C(\w_pixel_count[4] ), 
         .D(n36844), .Z(n4_adj_3975)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i1_4_lut_adj_515.init = 16'heccc;
    LUT4 i3_4_lut_adj_516 (.A(\w_pixel_count[0] ), .B(\w_pixel_count[1] ), 
         .C(\w_pixel_count[3] ), .D(\w_pixel_count[2] ), .Z(n36844)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut_adj_516.init = 16'hfffe;
    CCU2D pixel_count_19667_19668_add_4_11 (.A0(\w_pixel_count[9] ), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(\w_pixel_count[10] ), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n36657), .S0(n49[9]), .S1(n49[10]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam pixel_count_19667_19668_add_4_11.INIT0 = 16'hfaaa;
    defparam pixel_count_19667_19668_add_4_11.INIT1 = 16'hfaaa;
    defparam pixel_count_19667_19668_add_4_11.INJECT1_0 = "NO";
    defparam pixel_count_19667_19668_add_4_11.INJECT1_1 = "NO";
    CCU2D pixel_count_19667_19668_add_4_9 (.A0(\w_pixel_count[7] ), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(\w_pixel_count[8] ), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n36656), .COUT(n36657), .S0(n49[7]), 
          .S1(n49[8]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam pixel_count_19667_19668_add_4_9.INIT0 = 16'hfaaa;
    defparam pixel_count_19667_19668_add_4_9.INIT1 = 16'hfaaa;
    defparam pixel_count_19667_19668_add_4_9.INJECT1_0 = "NO";
    defparam pixel_count_19667_19668_add_4_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_317_3_lut_4_lut (.A(n41523), .B(w_line_count_c[9]), 
         .C(w_line_count[7]), .D(w_line_count_c[8]), .Z(n41404)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_317_3_lut_4_lut.init = 16'hfffe;
    LUT4 i29991_4_lut_4_lut (.A(n41523), .B(w_line_count_c[9]), .C(n38869), 
         .D(w_line_count_c[8]), .Z(n32575)) /* synthesis lut_function=(A+(B (C+(D)))) */ ;
    defparam i29991_4_lut_4_lut.init = 16'heeea;
    CCU2D pixel_count_19667_19668_add_4_7 (.A0(\w_pixel_count[5] ), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(\w_pixel_count[6] ), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n36655), .COUT(n36656), .S0(n49[5]), 
          .S1(n49[6]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam pixel_count_19667_19668_add_4_7.INIT0 = 16'hfaaa;
    defparam pixel_count_19667_19668_add_4_7.INIT1 = 16'hfaaa;
    defparam pixel_count_19667_19668_add_4_7.INJECT1_0 = "NO";
    defparam pixel_count_19667_19668_add_4_7.INJECT1_1 = "NO";
    CCU2D pixel_count_19667_19668_add_4_5 (.A0(\w_pixel_count[3] ), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(\w_pixel_count[4] ), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n36654), .COUT(n36655), .S0(n49[3]), 
          .S1(n49[4]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam pixel_count_19667_19668_add_4_5.INIT0 = 16'hfaaa;
    defparam pixel_count_19667_19668_add_4_5.INIT1 = 16'hfaaa;
    defparam pixel_count_19667_19668_add_4_5.INJECT1_0 = "NO";
    defparam pixel_count_19667_19668_add_4_5.INJECT1_1 = "NO";
    LUT4 i29935_3_lut_4_lut (.A(n41521), .B(w_line_count[4]), .C(\w_line_count[5] ), 
         .D(n41522), .Z(n32519)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;
    defparam i29935_3_lut_4_lut.init = 16'hf800;
    LUT4 i36647_3_lut_4_lut (.A(n41522), .B(n41520), .C(n41524), .D(w_line_count[2]), 
         .Z(n39197)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i36647_3_lut_4_lut.init = 16'h8880;
    LUT4 i27712_4_lut_4_lut (.A(n41522), .B(n41520), .C(\w_line_count[5] ), 
         .D(w_line_count[2]), .Z(n32466)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i27712_4_lut_4_lut.init = 16'ha8a0;
    CCU2D pixel_count_19667_19668_add_4_3 (.A0(\w_pixel_count[1] ), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(\w_pixel_count[2] ), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n36653), .COUT(n36654), .S0(n49[1]), 
          .S1(n49[2]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam pixel_count_19667_19668_add_4_3.INIT0 = 16'hfaaa;
    defparam pixel_count_19667_19668_add_4_3.INIT1 = 16'hfaaa;
    defparam pixel_count_19667_19668_add_4_3.INJECT1_0 = "NO";
    defparam pixel_count_19667_19668_add_4_3.INJECT1_1 = "NO";
    CCU2D pixel_count_19667_19668_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(\w_pixel_count[0] ), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n36653), .S1(n49[0]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/hvsync.v(42[19:37])
    defparam pixel_count_19667_19668_add_4_1.INIT0 = 16'hF000;
    defparam pixel_count_19667_19668_add_4_1.INIT1 = 16'h0555;
    defparam pixel_count_19667_19668_add_4_1.INJECT1_0 = "NO";
    defparam pixel_count_19667_19668_add_4_1.INJECT1_1 = "NO";
    PFUMX i38621 (.BLUT(n41615), .ALUT(n41616), .C0(\w_pixel_count[7] ), 
          .Z(n41617));
    
endmodule
//
// Verilog Description of module mico_cpu
//

module mico_cpu (\counter[2]_adj_101 , w_clk_cpu, reset_n_N_45, n41488, 
            sram_wen_N_3273, n42726, sramsram_data_in, sram_adr_c_0, 
            sramsram_data_out, sram_adr_c_18, sram_adr_c_17, sram_adr_c_16, 
            sram_adr_c_15, sram_adr_c_14, sram_adr_c_13, sram_adr_c_12, 
            sram_adr_c_11, sram_adr_c_10, sram_adr_c_9, sram_adr_c_8, 
            sram_adr_c_7, sram_adr_c_6, sram_adr_c_5, sram_adr_c_4, 
            sram_adr_c_3, sram_adr_c_2, sram_adr_c_1, sram_oen_c, \counter[0] , 
            \counter[1] , \counter[2] , \counter[4] , \counter[5] , 
            \counter[6] , \counter[7] , \counter[8] , \counter[9] , 
            \counter[10] , \counter[11] , \counter[12] , \counter[13] , 
            \counter[14] , \counter[15] , \counter[3] , GND_net, w_result, 
            read_idx_0_d, n23059, n23091, n23058, n23090, n23067, 
            n23099, n23068, n23100, n42734, n42738, read_idx_1_d, 
            n23069, n23101, n42732, n23070, n23102, n23071, n23103, 
            n23072, n23104, n41470, write_idx_w, n23185, n23186, 
            n23073, n23105, n23074, n23106, n23075, n23107, n23076, 
            n23108, n22885, reg_data_1, n23056, n23088, n23057, 
            n23089, n22999, n22877, n22874, n23053, n23085, n23054, 
            n23086, n23060, n23092, n23061, n23093, n23062, n23094, 
            n23063, n23095, n23064, n23096, n23065, n23097, n23066, 
            n23098, n23052, n23084, n23055, n23087, n23077, n23109, 
            n23078, n23110, n23079, n23111, n23080, n23112, n23081, 
            n23113, n23082, n23114, n23083, n23115, VCC_net) /* synthesis syn_module_defined=1 */ ;
    output \counter[2]_adj_101 ;
    input w_clk_cpu;
    input reset_n_N_45;
    output n41488;
    output sram_wen_N_3273;
    input n42726;
    input [7:0]sramsram_data_in;
    output sram_adr_c_0;
    output [7:0]sramsram_data_out;
    output sram_adr_c_18;
    output sram_adr_c_17;
    output sram_adr_c_16;
    output sram_adr_c_15;
    output sram_adr_c_14;
    output sram_adr_c_13;
    output sram_adr_c_12;
    output sram_adr_c_11;
    output sram_adr_c_10;
    output sram_adr_c_9;
    output sram_adr_c_8;
    output sram_adr_c_7;
    output sram_adr_c_6;
    output sram_adr_c_5;
    output sram_adr_c_4;
    output sram_adr_c_3;
    output sram_adr_c_2;
    output sram_adr_c_1;
    output sram_oen_c;
    output \counter[0] ;
    output \counter[1] ;
    output \counter[2] ;
    output \counter[4] ;
    output \counter[5] ;
    output \counter[6] ;
    output \counter[7] ;
    output \counter[8] ;
    output \counter[9] ;
    output \counter[10] ;
    output \counter[11] ;
    output \counter[12] ;
    output \counter[13] ;
    output \counter[14] ;
    output \counter[15] ;
    output \counter[3] ;
    input GND_net;
    output [31:0]w_result;
    output [4:0]read_idx_0_d;
    input n23059;
    input n23091;
    input n23058;
    input n23090;
    input n23067;
    input n23099;
    input n23068;
    input n23100;
    output n42734;
    output n42738;
    output [4:0]read_idx_1_d;
    input n23069;
    input n23101;
    output n42732;
    input n23070;
    input n23102;
    input n23071;
    input n23103;
    input n23072;
    input n23104;
    output n41470;
    output [4:0]write_idx_w;
    output n23185;
    output n23186;
    input n23073;
    input n23105;
    input n23074;
    input n23106;
    input n23075;
    input n23107;
    input n23076;
    input n23108;
    input n22885;
    input [31:0]reg_data_1;
    input n23056;
    input n23088;
    input n23057;
    input n23089;
    input n22999;
    output n22877;
    output n22874;
    input n23053;
    input n23085;
    input n23054;
    input n23086;
    input n23060;
    input n23092;
    input n23061;
    input n23093;
    input n23062;
    input n23094;
    input n23063;
    input n23095;
    input n23064;
    input n23096;
    input n23065;
    input n23097;
    input n23066;
    input n23098;
    input n23052;
    input n23084;
    input n23055;
    input n23087;
    input n23077;
    input n23109;
    input n23078;
    input n23110;
    input n23079;
    input n23111;
    input n23080;
    input n23112;
    input n23081;
    input n23113;
    input n23082;
    input n23114;
    input n23083;
    input n23115;
    input VCC_net;
    
    wire w_clk_cpu /* synthesis SET_AS_NETWORK=w_clk_cpu, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(22[6:15])
    
    wire n41442;
    wire [31:0]SHAREDBUS_ADR_I;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(348[13:28])
    
    wire n21, LM32I_CYC_O, n38871, n41479;
    wire [0:0]n76;
    
    wire i_cyc_o_N_1759;
    wire [31:0]sramASRAM_DAT_O;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(396[13:28])
    
    wire n41398, n38745, n38731, n38733, n38747;
    wire [0:0]n4;
    
    wire n41362, n7, n41501, n41353, n38735, n38757, n38737, n41393, 
        n41453, sram_data_out_nxt_7__N_3203, n38749, n38739, n38755, 
        n38741, n38751, n38743, n22, n38759, n38729, n38730, n38732, 
        n38734, n38736, n38738, n38740, n38742, n38744, n38746, 
        n38748, n38750, n38752, n38754, n14, n38756, n38758, n38760, 
        n38753, n41366, n38717, n41385;
    wire [2:0]n30;
    wire [2:0]n5;
    
    wire counter_2__N_178, n41370, n35, LM32DEBUG_ACK_O;
    wire [31:0]SHAREDBUS_ACK_O_N_81;
    
    wire n41421, gpioGPIO_ACK_O, n7_adj_3941;
    wire [31:0]SHAREDBUS_DAT_O;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(350[13:28])
    
    wire n7_adj_3942, n7_adj_3943, n7_adj_3944, n7_adj_3945, n7_adj_3946, 
        n7_adj_3947, n7_adj_3948, n7_adj_3949, n7_adj_3950, n7_adj_3951, 
        n7_adj_3952, n7_adj_3953, n7_adj_3954, n7_adj_3955, n7_adj_3956, 
        n7_adj_3957, n7_adj_3958, n7_adj_3959, n7_adj_3960, n7_adj_3961, 
        n39983, n17, n7_adj_3962, n16, n7_adj_3963, n7_adj_3964, 
        n7_adj_3965, n7_adj_3966, n7_adj_3967, n7_adj_3968, n7_adj_3969, 
        n7_adj_3970, n7_adj_3971, n41422, state_nxt_1__N_3154, n41356, 
        n7_adj_3972;
    wire [0:0]n1;
    
    wire n41352, n40733, n40734, n42723, n183, LM32D_CYC_O, n41490, 
        data_bus_error_exception_N_1225, wb_load_complete_N_2129, n41435, 
        n23, n10;
    wire [15:0]n21518;
    
    wire n41405, n7_adj_3973, n36822;
    wire [3:0]SHAREDBUS_SEL_I;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(351[12:27])
    
    wire n41344, tmp_ack_o, n24342, n28684, \genblk5.tmp_ack_o_d , 
        w_clk_cpu_enable_900, n26128;
    wire [31:0]LM32D_ADR_O;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(376[13:24])
    
    wire n41412;
    wire [3:0]LM32D_SEL_O;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(379[12:23])
    wire [1:0]selected;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(244[15:23])
    
    wire n41424, n38761, PIO_OUT_7__N_3327, n41423, n25515, n25664, 
        w_clk_cpu_enable_303, n41363, n24709, n39016;
    wire [31:0]LM32D_DAT_O;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(377[13:24])
    
    wire n36688, n22230, n38998, n31536, n37005, n39018, n41429, 
        n41390, n41392, n41469, n41455;
    wire [31:0]data;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(105[23:27])
    wire [31:0]SHAREDBUS_DAT_I;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(349[13:28])
    wire [7:0]n96;
    wire [31:0]tmp_dat_o_nxt_31__N_3207;
    
    wire LM32D_WE_O, n41426, PIO_OUT_15__N_3318;
    wire [1:0]selected_1__N_344;
    wire [31:0]LM32I_ADR_O;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(363[13:24])
    
    wire LM32D_STB_O;
    wire [7:0]n87;
    
    wire bus_error_f_N_1764;
    
    LUT4 i8_4_lut (.A(n41442), .B(SHAREDBUS_ADR_I[12]), .C(SHAREDBUS_ADR_I[8]), 
         .D(SHAREDBUS_ADR_I[5]), .Z(n21)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(567[23:68])
    defparam i8_4_lut.init = 16'hfffd;
    LUT4 i29503_3_lut_4_lut (.A(LM32I_CYC_O), .B(n38871), .C(n41479), 
         .D(n76[0]), .Z(i_cyc_o_N_1759)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i29503_3_lut_4_lut.init = 16'hf080;
    LUT4 i1_2_lut_4_lut_4_lut (.A(n41442), .B(sramASRAM_DAT_O[5]), .C(SHAREDBUS_ADR_I[20]), 
         .D(n41398), .Z(n38745)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_444 (.A(n41442), .B(sramASRAM_DAT_O[6]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38731)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_444.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_445 (.A(n41442), .B(sramASRAM_DAT_O[7]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38733)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_445.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_446 (.A(n41442), .B(sramASRAM_DAT_O[8]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38747)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_446.init = 16'h0004;
    LUT4 sram_addr_nxt_18__N_3070_I_0_3_lut_rep_266_4_lut (.A(n4[0]), .B(n41362), 
         .C(n7), .D(n41501), .Z(n41353)) /* synthesis lut_function=(!(A (B (C (D))+!B (D))+!A (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(590[14:44])
    defparam sram_addr_nxt_18__N_3070_I_0_3_lut_rep_266_4_lut.init = 16'h08ff;
    LUT4 i1_2_lut_4_lut_4_lut_adj_447 (.A(n41442), .B(sramASRAM_DAT_O[9]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38735)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_447.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_448 (.A(n41442), .B(sramASRAM_DAT_O[11]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38757)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_448.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_449 (.A(n41442), .B(sramASRAM_DAT_O[12]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38737)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_449.init = 16'h0004;
    LUT4 i2_3_lut_4_lut (.A(n4[0]), .B(n41362), .C(n41393), .D(n41453), 
         .Z(sram_data_out_nxt_7__N_3203)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(590[14:44])
    defparam i2_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_4_lut_4_lut_adj_450 (.A(n41442), .B(sramASRAM_DAT_O[13]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38749)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_450.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_451 (.A(n41442), .B(sramASRAM_DAT_O[14]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38739)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_451.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_452 (.A(n41442), .B(sramASRAM_DAT_O[15]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38755)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_452.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_453 (.A(n41442), .B(sramASRAM_DAT_O[16]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38741)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_453.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_454 (.A(n41442), .B(sramASRAM_DAT_O[17]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38751)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_454.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_455 (.A(n41442), .B(sramASRAM_DAT_O[18]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38743)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_455.init = 16'h0004;
    LUT4 i9_4_lut (.A(SHAREDBUS_ADR_I[4]), .B(SHAREDBUS_ADR_I[6]), .C(SHAREDBUS_ADR_I[20]), 
         .D(SHAREDBUS_ADR_I[9]), .Z(n22)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(567[23:68])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_4_lut_adj_456 (.A(n41442), .B(sramASRAM_DAT_O[19]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38759)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_456.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_457 (.A(n41442), .B(sramASRAM_DAT_O[20]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38729)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_457.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_458 (.A(n41442), .B(sramASRAM_DAT_O[21]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38730)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_458.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_459 (.A(n41442), .B(sramASRAM_DAT_O[22]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38732)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_459.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_460 (.A(n41442), .B(sramASRAM_DAT_O[23]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38734)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_460.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_461 (.A(n41442), .B(sramASRAM_DAT_O[24]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38736)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_461.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_462 (.A(n41442), .B(sramASRAM_DAT_O[25]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38738)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_462.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_463 (.A(n41442), .B(sramASRAM_DAT_O[26]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38740)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_463.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_464 (.A(n41442), .B(sramASRAM_DAT_O[27]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38742)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_464.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_465 (.A(n41442), .B(sramASRAM_DAT_O[29]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38744)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_465.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_466 (.A(n41442), .B(sramASRAM_DAT_O[30]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38746)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_466.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_467 (.A(n41442), .B(sramASRAM_DAT_O[31]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38748)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_467.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_468 (.A(n41442), .B(sramASRAM_DAT_O[28]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38750)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_468.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_469 (.A(n41442), .B(sramASRAM_DAT_O[10]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38752)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_469.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_470 (.A(n41442), .B(sramASRAM_DAT_O[4]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38754)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_470.init = 16'h0004;
    LUT4 i1_2_lut (.A(SHAREDBUS_ADR_I[10]), .B(SHAREDBUS_ADR_I[7]), .Z(n14)) /* synthesis lut_function=(A+(B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(567[23:68])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i1_2_lut_4_lut_4_lut_adj_471 (.A(n41442), .B(sramASRAM_DAT_O[1]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38756)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_471.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_472 (.A(n41442), .B(sramASRAM_DAT_O[0]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38758)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_472.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_473 (.A(n41442), .B(sramASRAM_DAT_O[2]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38760)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_473.init = 16'h0004;
    LUT4 i1_2_lut_4_lut_4_lut_adj_474 (.A(n41442), .B(sramASRAM_DAT_O[3]), 
         .C(SHAREDBUS_ADR_I[20]), .D(n41398), .Z(n38753)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_474.init = 16'h0004;
    LUT4 i1_4_lut_4_lut (.A(n41366), .B(n38717), .C(SHAREDBUS_ADR_I[20]), 
         .D(n41385), .Z(n38871)) /* synthesis lut_function=(!(A+!(B (C+(D))+!B (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(605[22:82])
    defparam i1_4_lut_4_lut.init = 16'h5540;
    LUT4 i34116_3_lut (.A(\counter[2]_adj_101 ), .B(n30[1]), .C(n30[0]), 
         .Z(n5[2])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(435[15:29])
    defparam i34116_3_lut.init = 16'h6a6a;
    LUT4 i34109_2_lut (.A(n30[1]), .B(n30[0]), .Z(n5[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(435[15:29])
    defparam i34109_2_lut.init = 16'h6666;
    LUT4 i34107_1_lut (.A(n30[0]), .Z(n5[0])) /* synthesis lut_function=(!(A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(435[15:29])
    defparam i34107_1_lut.init = 16'h5555;
    FD1P3DX counter_19665__i0 (.D(n5[0]), .SP(counter_2__N_178), .CK(w_clk_cpu), 
            .CD(reset_n_N_45), .Q(n30[0]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(435[15:29])
    defparam counter_19665__i0.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_298 (.A(n41398), .B(n41442), .Z(n41385)) /* synthesis lut_function=(A+(B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(567[23:68])
    defparam i1_2_lut_rep_298.init = 16'heeee;
    LUT4 i1_2_lut_rep_283_3_lut (.A(n41398), .B(n41442), .C(SHAREDBUS_ADR_I[20]), 
         .Z(n41370)) /* synthesis lut_function=(A+(B+(C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(567[23:68])
    defparam i1_2_lut_rep_283_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut (.A(n38717), .B(n41398), .C(n41442), .D(SHAREDBUS_ADR_I[20]), 
         .Z(n35)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(567[23:68])
    defparam i1_4_lut.init = 16'hfeff;
    PFUMX mux_6_i1 (.BLUT(LM32DEBUG_ACK_O), .ALUT(SHAREDBUS_ACK_O_N_81[0]), 
          .C0(n35), .Z(n76[0])) /* synthesis LSE_LINE_FILE_ID=7, LSE_LCOL=10, LSE_RCOL=2, LSE_LLINE=34, LSE_RLINE=44 */ ;
    LUT4 mux_83_i1_4_lut (.A(n41421), .B(gpioGPIO_ACK_O), .C(n41370), 
         .D(n41366), .Z(SHAREDBUS_ACK_O_N_81[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(505[1] 507[2])
    defparam mux_83_i1_4_lut.init = 16'hca0a;
    PFUMX i15 (.BLUT(n7_adj_3941), .ALUT(n38753), .C0(n35), .Z(SHAREDBUS_DAT_O[3]));
    PFUMX i15_adj_475 (.BLUT(n7_adj_3942), .ALUT(n38760), .C0(n35), .Z(SHAREDBUS_DAT_O[2]));
    PFUMX i15_adj_476 (.BLUT(n7_adj_3943), .ALUT(n38758), .C0(n35), .Z(SHAREDBUS_DAT_O[0]));
    PFUMX i15_adj_477 (.BLUT(n7_adj_3944), .ALUT(n38756), .C0(n35), .Z(SHAREDBUS_DAT_O[1]));
    PFUMX i15_adj_478 (.BLUT(n7_adj_3945), .ALUT(n38754), .C0(n35), .Z(SHAREDBUS_DAT_O[4]));
    PFUMX i15_adj_479 (.BLUT(n7_adj_3946), .ALUT(n38752), .C0(n35), .Z(SHAREDBUS_DAT_O[10]));
    PFUMX i15_adj_480 (.BLUT(n7_adj_3947), .ALUT(n38750), .C0(n35), .Z(SHAREDBUS_DAT_O[28]));
    PFUMX i15_adj_481 (.BLUT(n7_adj_3948), .ALUT(n38748), .C0(n35), .Z(SHAREDBUS_DAT_O[31]));
    PFUMX i15_adj_482 (.BLUT(n7_adj_3949), .ALUT(n38746), .C0(n35), .Z(SHAREDBUS_DAT_O[30]));
    PFUMX i15_adj_483 (.BLUT(n7_adj_3950), .ALUT(n38744), .C0(n35), .Z(SHAREDBUS_DAT_O[29]));
    PFUMX i15_adj_484 (.BLUT(n7_adj_3951), .ALUT(n38742), .C0(n35), .Z(SHAREDBUS_DAT_O[27]));
    PFUMX i15_adj_485 (.BLUT(n7_adj_3952), .ALUT(n38740), .C0(n35), .Z(SHAREDBUS_DAT_O[26]));
    PFUMX i15_adj_486 (.BLUT(n7_adj_3953), .ALUT(n38738), .C0(n35), .Z(SHAREDBUS_DAT_O[25]));
    PFUMX i15_adj_487 (.BLUT(n7_adj_3954), .ALUT(n38736), .C0(n35), .Z(SHAREDBUS_DAT_O[24]));
    PFUMX i15_adj_488 (.BLUT(n7_adj_3955), .ALUT(n38734), .C0(n35), .Z(SHAREDBUS_DAT_O[23]));
    PFUMX i15_adj_489 (.BLUT(n7_adj_3956), .ALUT(n38732), .C0(n35), .Z(SHAREDBUS_DAT_O[22]));
    PFUMX i15_adj_490 (.BLUT(n7_adj_3957), .ALUT(n38730), .C0(n35), .Z(SHAREDBUS_DAT_O[21]));
    PFUMX i15_adj_491 (.BLUT(n7_adj_3958), .ALUT(n38729), .C0(n35), .Z(SHAREDBUS_DAT_O[20]));
    PFUMX i15_adj_492 (.BLUT(n7_adj_3959), .ALUT(n38759), .C0(n35), .Z(SHAREDBUS_DAT_O[19]));
    PFUMX i15_adj_493 (.BLUT(n7_adj_3960), .ALUT(n38743), .C0(n35), .Z(SHAREDBUS_DAT_O[18]));
    PFUMX i15_adj_494 (.BLUT(n7_adj_3961), .ALUT(n38751), .C0(n35), .Z(SHAREDBUS_DAT_O[17]));
    LUT4 i37902_3_lut_4_lut (.A(SHAREDBUS_ADR_I[20]), .B(n41385), .C(n41488), 
         .D(n39983), .Z(sram_wen_N_3273)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(567[23:68])
    defparam i37902_3_lut_4_lut.init = 16'hfffe;
    LUT4 counter_2__I_0_1_lut (.A(\counter[2]_adj_101 ), .Z(counter_2__N_178)) /* synthesis lut_function=(!(A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(429[18:29])
    defparam counter_2__I_0_1_lut.init = 16'h5555;
    LUT4 i7_4_lut (.A(SHAREDBUS_ADR_I[23]), .B(SHAREDBUS_ADR_I[29]), .C(SHAREDBUS_ADR_I[28]), 
         .D(SHAREDBUS_ADR_I[27]), .Z(n17)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i7_4_lut.init = 16'hfffe;
    PFUMX i15_adj_495 (.BLUT(n7_adj_3962), .ALUT(n38741), .C0(n35), .Z(SHAREDBUS_DAT_O[16]));
    LUT4 i6_4_lut (.A(SHAREDBUS_ADR_I[24]), .B(SHAREDBUS_ADR_I[25]), .C(SHAREDBUS_ADR_I[26]), 
         .D(SHAREDBUS_ADR_I[22]), .Z(n16)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i6_4_lut.init = 16'hfffe;
    PFUMX i15_adj_496 (.BLUT(n7_adj_3963), .ALUT(n38755), .C0(n35), .Z(SHAREDBUS_DAT_O[15]));
    LUT4 i9_4_lut_rep_311 (.A(n17), .B(SHAREDBUS_ADR_I[21]), .C(n16), 
         .D(SHAREDBUS_ADR_I[30]), .Z(n41398)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i9_4_lut_rep_311.init = 16'hfffe;
    PFUMX i15_adj_497 (.BLUT(n7_adj_3964), .ALUT(n38739), .C0(n35), .Z(SHAREDBUS_DAT_O[14]));
    PFUMX i15_adj_498 (.BLUT(n7_adj_3965), .ALUT(n38749), .C0(n35), .Z(SHAREDBUS_DAT_O[13]));
    PFUMX i15_adj_499 (.BLUT(n7_adj_3966), .ALUT(n38737), .C0(n35), .Z(SHAREDBUS_DAT_O[12]));
    PFUMX i15_adj_500 (.BLUT(n7_adj_3967), .ALUT(n38757), .C0(n35), .Z(SHAREDBUS_DAT_O[11]));
    PFUMX i15_adj_501 (.BLUT(n7_adj_3968), .ALUT(n38735), .C0(n35), .Z(SHAREDBUS_DAT_O[9]));
    PFUMX i15_adj_502 (.BLUT(n7_adj_3969), .ALUT(n38747), .C0(n35), .Z(SHAREDBUS_DAT_O[8]));
    PFUMX i15_adj_503 (.BLUT(n7_adj_3970), .ALUT(n38733), .C0(n35), .Z(SHAREDBUS_DAT_O[7]));
    PFUMX i15_adj_504 (.BLUT(n7_adj_3971), .ALUT(n38731), .C0(n35), .Z(SHAREDBUS_DAT_O[6]));
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n41421), .B(n41422), .C(n41385), 
         .D(SHAREDBUS_ADR_I[20]), .Z(state_nxt_1__N_3154)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h0004;
    LUT4 i1_2_lut_rep_269_3_lut_4_lut_4_lut (.A(n41421), .B(n4[0]), .C(n41385), 
         .D(SHAREDBUS_ADR_I[20]), .Z(n41356)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i1_2_lut_rep_269_3_lut_4_lut_4_lut.init = 16'h0004;
    PFUMX i15_adj_505 (.BLUT(n7_adj_3972), .ALUT(n38745), .C0(n35), .Z(SHAREDBUS_DAT_O[5]));
    LUT4 i1_2_lut_rep_265 (.A(n1[0]), .B(n38871), .Z(n41352)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_265.init = 16'h8888;
    FD1P3DX counter_19665__i2 (.D(n42726), .SP(n5[2]), .CK(w_clk_cpu), 
            .CD(reset_n_N_45), .Q(\counter[2]_adj_101 ));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(435[15:29])
    defparam counter_19665__i2.GSR = "DISABLED";
    FD1P3DX counter_19665__i1 (.D(n5[1]), .SP(counter_2__N_178), .CK(w_clk_cpu), 
            .CD(reset_n_N_45), .Q(n30[1]));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(435[15:29])
    defparam counter_19665__i1.GSR = "DISABLED";
    LUT4 b_c_bdd_2_lut_38237_3_lut_4_lut_4_lut (.A(n41421), .B(n4[0]), .C(n40733), 
         .D(n41370), .Z(n40734)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam b_c_bdd_2_lut_38237_3_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i119_2_lut_3_lut_4_lut_4_lut (.A(n41421), .B(n4[0]), .C(n42723), 
         .D(n41370), .Z(n183)) /* synthesis lut_function=(!(A (C)+!A (B (C+!(D))+!B (C)))) */ ;
    defparam i119_2_lut_3_lut_4_lut_4_lut.init = 16'h0f0b;
    LUT4 i2_3_lut_4_lut_adj_506 (.A(n1[0]), .B(n38871), .C(LM32D_CYC_O), 
         .D(n41490), .Z(data_bus_error_exception_N_1225)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i2_3_lut_4_lut_adj_506.init = 16'h0080;
    LUT4 i37913_2_lut_rep_275_3_lut_4_lut_4_lut (.A(n41421), .B(SHAREDBUS_ADR_I[20]), 
         .C(n41442), .D(n41398), .Z(n41362)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i37913_2_lut_rep_275_3_lut_4_lut_4_lut.init = 16'h0001;
    LUT4 i29464_3_lut_4_lut (.A(n1[0]), .B(n38871), .C(n41490), .D(n76[0]), 
         .Z(wb_load_complete_N_2129)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (C+!(D)))) */ ;
    defparam i29464_3_lut_4_lut.init = 16'h0f08;
    LUT4 i10_4_lut (.A(SHAREDBUS_ADR_I[11]), .B(n38717), .C(n41435), .D(n14), 
         .Z(n23)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(567[23:68])
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i5_3_lut (.A(SHAREDBUS_ADR_I[19]), .B(n10), .C(SHAREDBUS_ADR_I[17]), 
         .Z(n38717)) /* synthesis lut_function=(A+(B+(C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(567[23:68])
    defparam i5_3_lut.init = 16'hfefe;
    LUT4 i4_4_lut (.A(SHAREDBUS_ADR_I[14]), .B(SHAREDBUS_ADR_I[15]), .C(SHAREDBUS_ADR_I[18]), 
         .D(SHAREDBUS_ADR_I[16]), .Z(n10)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(567[23:68])
    defparam i4_4_lut.init = 16'hfffe;
    LUT4 i38050_4_lut_rep_279_4_lut (.A(n41398), .B(n22), .C(n21), .D(n23), 
         .Z(n41366)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(605[22:82])
    defparam i38050_4_lut_rep_279_4_lut.init = 16'h0001;
    \asram_top(SRAM_DATA_WIDTH=8,SRAM_ADDR_WIDTH=19,SRAM_BE_WIDTH=1,READ_LATENCY=2,WRITE_LATENCY=2,DATA_OUTPUT_REG=1)  sramASRAM_DAT_O_31__I_0 (.sramASRAM_DAT_O({sramASRAM_DAT_O}), 
            .sramsram_data_in({sramsram_data_in}), .n21531(n21518[3]), .n41405(n41405), 
            .n7(n7_adj_3973), .n41393(n41393), .n36822(n36822), .n41501(n41501), 
            .n7_adj_100(n7), .n41356(n41356), .\SHAREDBUS_SEL_I[1] (SHAREDBUS_SEL_I[1]), 
            .n41344(n41344), .w_clk_cpu(w_clk_cpu), .tmp_ack_o(tmp_ack_o), 
            .n41488(n41488), .n24342(n24342), .n28684(n28684), .sram_adr_c_0(sram_adr_c_0), 
            .\genblk5.tmp_ack_o_d (\genblk5.tmp_ack_o_d ), .n42723(n42723), 
            .sramsram_data_out({sramsram_data_out}), .w_clk_cpu_enable_900(w_clk_cpu_enable_900), 
            .n26128(n26128), .sram_adr_c_18(sram_adr_c_18), .\SHAREDBUS_ADR_I[18] (SHAREDBUS_ADR_I[18]), 
            .sram_adr_c_17(sram_adr_c_17), .\SHAREDBUS_ADR_I[17] (SHAREDBUS_ADR_I[17]), 
            .sram_adr_c_16(sram_adr_c_16), .\SHAREDBUS_ADR_I[16] (SHAREDBUS_ADR_I[16]), 
            .sram_adr_c_15(sram_adr_c_15), .\SHAREDBUS_ADR_I[15] (SHAREDBUS_ADR_I[15]), 
            .\SHAREDBUS_ADR_I[0] (SHAREDBUS_ADR_I[0]), .sram_adr_c_14(sram_adr_c_14), 
            .\SHAREDBUS_ADR_I[14] (SHAREDBUS_ADR_I[14]), .sram_adr_c_13(sram_adr_c_13), 
            .n41435(n41435), .\LM32D_ADR_O[1] (LM32D_ADR_O[1]), .n41412(n41412), 
            .sram_adr_c_12(sram_adr_c_12), .\SHAREDBUS_ADR_I[12] (SHAREDBUS_ADR_I[12]), 
            .sram_adr_c_11(sram_adr_c_11), .\SHAREDBUS_ADR_I[11] (SHAREDBUS_ADR_I[11]), 
            .sram_adr_c_10(sram_adr_c_10), .\SHAREDBUS_ADR_I[10] (SHAREDBUS_ADR_I[10]), 
            .sram_adr_c_9(sram_adr_c_9), .\SHAREDBUS_ADR_I[9] (SHAREDBUS_ADR_I[9]), 
            .n41353(n41353), .sram_adr_c_8(sram_adr_c_8), .\SHAREDBUS_ADR_I[8] (SHAREDBUS_ADR_I[8]), 
            .sram_adr_c_7(sram_adr_c_7), .\SHAREDBUS_ADR_I[7] (SHAREDBUS_ADR_I[7]), 
            .sram_adr_c_6(sram_adr_c_6), .\SHAREDBUS_ADR_I[6] (SHAREDBUS_ADR_I[6]), 
            .sram_adr_c_5(sram_adr_c_5), .\SHAREDBUS_ADR_I[5] (SHAREDBUS_ADR_I[5]), 
            .sram_adr_c_4(sram_adr_c_4), .\SHAREDBUS_ADR_I[4] (SHAREDBUS_ADR_I[4]), 
            .sram_adr_c_3(sram_adr_c_3), .\SHAREDBUS_ADR_I[3] (SHAREDBUS_ADR_I[3]), 
            .sram_adr_c_2(sram_adr_c_2), .\SHAREDBUS_ADR_I[2] (SHAREDBUS_ADR_I[2]), 
            .sram_adr_c_1(sram_adr_c_1), .LM32D_SEL_O({LM32D_SEL_O}), .selected({selected}), 
            .n41424(n41424), .n38761(n38761), .PIO_OUT_7__N_3327(PIO_OUT_7__N_3327), 
            .n41423(n41423), .n41490(n41490), .n25515(n25515), .n25664(n25664), 
            .w_clk_cpu_enable_303(w_clk_cpu_enable_303), .n41363(n41363), 
            .n24709(n24709), .n39016(n39016), .LM32D_DAT_O({LM32D_DAT_O}), 
            .n36688(n36688), .n183(n183), .n22230(n22230), .n38998(n38998), 
            .n31536(n31536), .sram_data_out_nxt_7__N_3203(sram_data_out_nxt_7__N_3203), 
            .n37005(n37005), .n39018(n39018), .n40734(n40734), .state_nxt_1__N_3154(state_nxt_1__N_3154), 
            .n41429(n41429), .n41390(n41390), .n40733(n40733), .n41453(n41453), 
            .n41392(n41392), .n41479(n41479), .n41469(n41469), .n41455(n41455), 
            .\data[28] (data[28]), .\SHAREDBUS_DAT_I[28] (SHAREDBUS_DAT_I[28]), 
            .n96({n96}), .\data[29] (data[29]), .\SHAREDBUS_DAT_I[29] (SHAREDBUS_DAT_I[29]), 
            .\data[30] (data[30]), .\SHAREDBUS_DAT_I[30] (SHAREDBUS_DAT_I[30]), 
            .\data[31] (data[31]), .\SHAREDBUS_DAT_I[31] (SHAREDBUS_DAT_I[31]), 
            .\data[27] (data[27]), .\SHAREDBUS_DAT_I[27] (SHAREDBUS_DAT_I[27]), 
            .\data[26] (data[26]), .\SHAREDBUS_DAT_I[26] (SHAREDBUS_DAT_I[26]), 
            .\data[25] (data[25]), .\SHAREDBUS_DAT_I[25] (SHAREDBUS_DAT_I[25]), 
            .\data[24] (data[24]), .\SHAREDBUS_DAT_I[24] (SHAREDBUS_DAT_I[24]), 
            .\tmp_dat_o_nxt_31__N_3207[19] (tmp_dat_o_nxt_31__N_3207[19]), 
            .LM32D_WE_O(LM32D_WE_O), .sram_oen_c(sram_oen_c), .n41426(n41426)) /* synthesis syn_module_defined=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(577[2] 598[36])
    \gpio(DATA_WIDTH=32'b0100000,INPUT_WIDTH=32'b01,OUTPUT_WIDTH=32'b01,EDGE=1,POSE_EDGE_IRQ=1,INPUT_PORTS_ONLY=0,OUTPUT_PORTS_ONLY=1)  gpioGPIO_DAT_O_31__I_0 (.gpioGPIO_ACK_O(gpioGPIO_ACK_O), 
            .n93({n4}), .n41366(n41366), .w_clk_cpu(w_clk_cpu), .\counter[0] (\counter[0] ), 
            .PIO_OUT_7__N_3327(PIO_OUT_7__N_3327), .\SHAREDBUS_DAT_I[24] (SHAREDBUS_DAT_I[24]), 
            .\counter[1] (\counter[1] ), .\SHAREDBUS_DAT_I[25] (SHAREDBUS_DAT_I[25]), 
            .\counter[2] (\counter[2] ), .\SHAREDBUS_DAT_I[26] (SHAREDBUS_DAT_I[26]), 
            .w_clk_cpu_enable_303(w_clk_cpu_enable_303), .\SHAREDBUS_ADR_I[2] (SHAREDBUS_ADR_I[2]), 
            .\SHAREDBUS_ADR_I[3] (SHAREDBUS_ADR_I[3]), .n38761(n38761), 
            .\counter[4] (\counter[4] ), .\SHAREDBUS_DAT_I[28] (SHAREDBUS_DAT_I[28]), 
            .\counter[5] (\counter[5] ), .\SHAREDBUS_DAT_I[29] (SHAREDBUS_DAT_I[29]), 
            .\counter[6] (\counter[6] ), .\SHAREDBUS_DAT_I[30] (SHAREDBUS_DAT_I[30]), 
            .\counter[7] (\counter[7] ), .\SHAREDBUS_DAT_I[31] (SHAREDBUS_DAT_I[31]), 
            .\counter[8] (\counter[8] ), .PIO_OUT_15__N_3318(PIO_OUT_15__N_3318), 
            .\SHAREDBUS_DAT_I[16] (SHAREDBUS_DAT_I[16]), .\counter[9] (\counter[9] ), 
            .\SHAREDBUS_DAT_I[17] (SHAREDBUS_DAT_I[17]), .\counter[10] (\counter[10] ), 
            .\SHAREDBUS_DAT_I[18] (SHAREDBUS_DAT_I[18]), .\counter[11] (\counter[11] ), 
            .\SHAREDBUS_DAT_I[19] (SHAREDBUS_DAT_I[19]), .\counter[12] (\counter[12] ), 
            .\SHAREDBUS_DAT_I[20] (SHAREDBUS_DAT_I[20]), .\counter[13] (\counter[13] ), 
            .\SHAREDBUS_DAT_I[21] (SHAREDBUS_DAT_I[21]), .\counter[14] (\counter[14] ), 
            .\SHAREDBUS_DAT_I[22] (SHAREDBUS_DAT_I[22]), .\counter[15] (\counter[15] ), 
            .\SHAREDBUS_DAT_I[23] (SHAREDBUS_DAT_I[23]), .\counter[3] (\counter[3] ), 
            .\SHAREDBUS_DAT_I[27] (SHAREDBUS_DAT_I[27])) /* synthesis syn_module_defined=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(623[2] 639[34])
    arbiter2 arbiter (.n41426(n41426), .n41405(n41405), .n41424(n41424), 
            .n31536(n31536), .selected({selected}), .\selected_1__N_344[0] (selected_1__N_344[0]), 
            .w_clk_cpu(w_clk_cpu), .LM32D_SEL_O({LM32D_SEL_O}), .LM32D_WE_O(LM32D_WE_O), 
            .w_clk_cpu_enable_303(w_clk_cpu_enable_303), .n92({n1}), .n39983(n39983), 
            .\LM32I_ADR_O[11] (LM32I_ADR_O[11]), .\LM32D_ADR_O[11] (LM32D_ADR_O[11]), 
            .\SHAREDBUS_ADR_I[11] (SHAREDBUS_ADR_I[11]), .n25515(n25515), 
            .n41392(n41392), .n38761(n38761), .PIO_OUT_15__N_3318(PIO_OUT_15__N_3318), 
            .n41344(n41344), .n22230(n22230), .\LM32I_ADR_O[5] (LM32I_ADR_O[5]), 
            .\LM32D_ADR_O[5] (LM32D_ADR_O[5]), .\SHAREDBUS_ADR_I[5] (SHAREDBUS_ADR_I[5]), 
            .\LM32I_ADR_O[8] (LM32I_ADR_O[8]), .\LM32D_ADR_O[8] (LM32D_ADR_O[8]), 
            .\SHAREDBUS_ADR_I[8] (SHAREDBUS_ADR_I[8]), .\LM32I_ADR_O[12] (LM32I_ADR_O[12]), 
            .\LM32D_ADR_O[12] (LM32D_ADR_O[12]), .\SHAREDBUS_ADR_I[12] (SHAREDBUS_ADR_I[12]), 
            .w_clk_cpu_enable_900(w_clk_cpu_enable_900), .n26128(n26128), 
            .\LM32I_ADR_O[17] (LM32I_ADR_O[17]), .\LM32D_ADR_O[17] (LM32D_ADR_O[17]), 
            .\SHAREDBUS_ADR_I[17] (SHAREDBUS_ADR_I[17]), .\LM32I_ADR_O[16] (LM32I_ADR_O[16]), 
            .\LM32D_ADR_O[16] (LM32D_ADR_O[16]), .\SHAREDBUS_ADR_I[16] (SHAREDBUS_ADR_I[16]), 
            .\LM32I_ADR_O[18] (LM32I_ADR_O[18]), .\LM32D_ADR_O[18] (LM32D_ADR_O[18]), 
            .\SHAREDBUS_ADR_I[18] (SHAREDBUS_ADR_I[18]), .\LM32I_ADR_O[15] (LM32I_ADR_O[15]), 
            .\LM32D_ADR_O[15] (LM32D_ADR_O[15]), .\SHAREDBUS_ADR_I[15] (SHAREDBUS_ADR_I[15]), 
            .\LM32I_ADR_O[14] (LM32I_ADR_O[14]), .\LM32D_ADR_O[14] (LM32D_ADR_O[14]), 
            .\SHAREDBUS_ADR_I[14] (SHAREDBUS_ADR_I[14]), .\LM32D_DAT_O[24] (LM32D_DAT_O[24]), 
            .\SHAREDBUS_DAT_I[24] (SHAREDBUS_DAT_I[24]), .\LM32D_DAT_O[25] (LM32D_DAT_O[25]), 
            .\SHAREDBUS_DAT_I[25] (SHAREDBUS_DAT_I[25]), .\SHAREDBUS_SEL_I[1] (SHAREDBUS_SEL_I[1]), 
            .n41429(n41429), .\LM32I_ADR_O[19] (LM32I_ADR_O[19]), .\LM32D_ADR_O[19] (LM32D_ADR_O[19]), 
            .\SHAREDBUS_ADR_I[19] (SHAREDBUS_ADR_I[19]), .\LM32I_ADR_O[7] (LM32I_ADR_O[7]), 
            .\LM32D_ADR_O[7] (LM32D_ADR_O[7]), .\SHAREDBUS_ADR_I[7] (SHAREDBUS_ADR_I[7]), 
            .\LM32I_ADR_O[10] (LM32I_ADR_O[10]), .\LM32D_ADR_O[10] (LM32D_ADR_O[10]), 
            .\SHAREDBUS_ADR_I[10] (SHAREDBUS_ADR_I[10]), .\LM32I_ADR_O[9] (LM32I_ADR_O[9]), 
            .\LM32D_ADR_O[9] (LM32D_ADR_O[9]), .\SHAREDBUS_ADR_I[9] (SHAREDBUS_ADR_I[9]), 
            .\LM32I_ADR_O[6] (LM32I_ADR_O[6]), .\LM32D_ADR_O[6] (LM32D_ADR_O[6]), 
            .\SHAREDBUS_ADR_I[6] (SHAREDBUS_ADR_I[6]), .\LM32I_ADR_O[4] (LM32I_ADR_O[4]), 
            .\LM32D_ADR_O[4] (LM32D_ADR_O[4]), .\SHAREDBUS_ADR_I[4] (SHAREDBUS_ADR_I[4]), 
            .\LM32I_ADR_O[31] (LM32I_ADR_O[31]), .\LM32D_ADR_O[31] (LM32D_ADR_O[31]), 
            .n41442(n41442), .n41423(n41423), .\LM32I_ADR_O[13] (LM32I_ADR_O[13]), 
            .\LM32D_ADR_O[13] (LM32D_ADR_O[13]), .n41435(n41435), .\LM32I_ADR_O[22] (LM32I_ADR_O[22]), 
            .\LM32D_ADR_O[22] (LM32D_ADR_O[22]), .\SHAREDBUS_ADR_I[22] (SHAREDBUS_ADR_I[22]), 
            .\LM32I_ADR_O[26] (LM32I_ADR_O[26]), .\LM32D_ADR_O[26] (LM32D_ADR_O[26]), 
            .\SHAREDBUS_ADR_I[26] (SHAREDBUS_ADR_I[26]), .\LM32I_ADR_O[25] (LM32I_ADR_O[25]), 
            .\LM32D_ADR_O[25] (LM32D_ADR_O[25]), .\SHAREDBUS_ADR_I[25] (SHAREDBUS_ADR_I[25]), 
            .\LM32I_ADR_O[24] (LM32I_ADR_O[24]), .\LM32D_ADR_O[24] (LM32D_ADR_O[24]), 
            .\SHAREDBUS_ADR_I[24] (SHAREDBUS_ADR_I[24]), .\LM32I_ADR_O[27] (LM32I_ADR_O[27]), 
            .\LM32D_ADR_O[27] (LM32D_ADR_O[27]), .\SHAREDBUS_ADR_I[27] (SHAREDBUS_ADR_I[27]), 
            .\LM32I_ADR_O[28] (LM32I_ADR_O[28]), .\LM32D_ADR_O[28] (LM32D_ADR_O[28]), 
            .\SHAREDBUS_ADR_I[28] (SHAREDBUS_ADR_I[28]), .\LM32D_DAT_O[26] (LM32D_DAT_O[26]), 
            .\SHAREDBUS_DAT_I[26] (SHAREDBUS_DAT_I[26]), .\LM32D_DAT_O[28] (LM32D_DAT_O[28]), 
            .\SHAREDBUS_DAT_I[28] (SHAREDBUS_DAT_I[28]), .\LM32I_ADR_O[29] (LM32I_ADR_O[29]), 
            .\LM32D_ADR_O[29] (LM32D_ADR_O[29]), .\SHAREDBUS_ADR_I[29] (SHAREDBUS_ADR_I[29]), 
            .\LM32D_DAT_O[29] (LM32D_DAT_O[29]), .\SHAREDBUS_DAT_I[29] (SHAREDBUS_DAT_I[29]), 
            .\LM32D_DAT_O[30] (LM32D_DAT_O[30]), .\SHAREDBUS_DAT_I[30] (SHAREDBUS_DAT_I[30]), 
            .\LM32D_DAT_O[31] (LM32D_DAT_O[31]), .\SHAREDBUS_DAT_I[31] (SHAREDBUS_DAT_I[31]), 
            .\LM32D_DAT_O[18] (LM32D_DAT_O[18]), .\SHAREDBUS_DAT_I[18] (SHAREDBUS_DAT_I[18]), 
            .\LM32D_DAT_O[19] (LM32D_DAT_O[19]), .\SHAREDBUS_DAT_I[19] (SHAREDBUS_DAT_I[19]), 
            .\LM32I_ADR_O[23] (LM32I_ADR_O[23]), .\LM32D_ADR_O[23] (LM32D_ADR_O[23]), 
            .\SHAREDBUS_ADR_I[23] (SHAREDBUS_ADR_I[23]), .\LM32I_ADR_O[30] (LM32I_ADR_O[30]), 
            .\LM32D_ADR_O[30] (LM32D_ADR_O[30]), .\SHAREDBUS_ADR_I[30] (SHAREDBUS_ADR_I[30]), 
            .\LM32D_DAT_O[20] (LM32D_DAT_O[20]), .\SHAREDBUS_DAT_I[20] (SHAREDBUS_DAT_I[20]), 
            .\LM32I_ADR_O[21] (LM32I_ADR_O[21]), .\LM32D_ADR_O[21] (LM32D_ADR_O[21]), 
            .\SHAREDBUS_ADR_I[21] (SHAREDBUS_ADR_I[21]), .\LM32I_ADR_O[2] (LM32I_ADR_O[2]), 
            .\LM32D_ADR_O[2] (LM32D_ADR_O[2]), .\SHAREDBUS_ADR_I[2] (SHAREDBUS_ADR_I[2]), 
            .\LM32D_DAT_O[21] (LM32D_DAT_O[21]), .\SHAREDBUS_DAT_I[21] (SHAREDBUS_DAT_I[21]), 
            .\LM32I_ADR_O[3] (LM32I_ADR_O[3]), .\LM32D_ADR_O[3] (LM32D_ADR_O[3]), 
            .\SHAREDBUS_ADR_I[3] (SHAREDBUS_ADR_I[3]), .\LM32D_DAT_O[22] (LM32D_DAT_O[22]), 
            .\SHAREDBUS_DAT_I[22] (SHAREDBUS_DAT_I[22]), .\LM32D_DAT_O[23] (LM32D_DAT_O[23]), 
            .\SHAREDBUS_DAT_I[23] (SHAREDBUS_DAT_I[23]), .\LM32D_DAT_O[27] (LM32D_DAT_O[27]), 
            .\SHAREDBUS_DAT_I[27] (SHAREDBUS_DAT_I[27]), .\LM32I_ADR_O[20] (LM32I_ADR_O[20]), 
            .\LM32D_ADR_O[20] (LM32D_ADR_O[20]), .\SHAREDBUS_ADR_I[20] (SHAREDBUS_ADR_I[20]), 
            .LM32I_CYC_O(LM32I_CYC_O), .LM32D_CYC_O(LM32D_CYC_O), .LM32D_STB_O(LM32D_STB_O), 
            .n93({n4}), .n41479(n41479), .n38998(n38998), .n41393(n41393), 
            .n41469(n41469), .\data[19] (data[19]), .n87({n87}), .n41390(n41390), 
            .n41363(n41363), .\SHAREDBUS_DAT_I[16] (SHAREDBUS_DAT_I[16]), 
            .\data[16] (data[16]), .\SHAREDBUS_DAT_I[17] (SHAREDBUS_DAT_I[17]), 
            .\data[17] (data[17]), .\data[23] (data[23]), .\data[18] (data[18]), 
            .\data[22] (data[22]), .\data[20] (data[20]), .\data[21] (data[21]), 
            .n41490(n41490), .n24709(n24709), .n41412(n41412), .n41455(n41455), 
            .\LM32D_DAT_O[17] (LM32D_DAT_O[17]), .tmp_ack_o(tmp_ack_o), 
            .\genblk5.tmp_ack_o_d (\genblk5.tmp_ack_o_d ), .n41421(n41421), 
            .n42723(n42723), .n25664(n25664), .n36688(n36688), .n24342(n24342), 
            .n36822(n36822), .n37005(n37005), .\LM32D_DAT_O[16] (LM32D_DAT_O[16]), 
            .n41352(n41352), .n76({n76}), .n39016(n39016), .n39018(n39018), 
            .n21531(n21518[3]), .\sramsram_data_in[3] (sramsram_data_in[3]), 
            .n7(n7_adj_3973), .n28684(n28684), .\tmp_dat_o_nxt_31__N_3207[19] (tmp_dat_o_nxt_31__N_3207[19]), 
            .n38871(n38871), .bus_error_f_N_1764(bus_error_f_N_1764), .\LM32D_ADR_O[0] (LM32D_ADR_O[0]), 
            .\SHAREDBUS_ADR_I[0] (SHAREDBUS_ADR_I[0])) /* synthesis syn_module_defined=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(451[1] 492[20])
    lm32_top LM32I_ADR_O_31__I_0 (.GND_net(GND_net), .n41435(n41435), .n7(n7_adj_3972), 
            .n7_adj_64(n7_adj_3971), .n7_adj_65(n7_adj_3970), .n7_adj_66(n7_adj_3969), 
            .n7_adj_67(n7_adj_3968), .n7_adj_68(n7_adj_3967), .n7_adj_69(n7_adj_3966), 
            .n7_adj_70(n7_adj_3965), .n7_adj_71(n7_adj_3964), .n7_adj_72(n7_adj_3963), 
            .n7_adj_73(n7_adj_3962), .n7_adj_74(n7_adj_3961), .n7_adj_75(n7_adj_3960), 
            .n7_adj_76(n7_adj_3959), .n7_adj_77(n7_adj_3958), .n7_adj_78(n7_adj_3957), 
            .n7_adj_79(n7_adj_3956), .n7_adj_80(n7_adj_3955), .n7_adj_81(n7_adj_3954), 
            .n7_adj_82(n7_adj_3953), .n7_adj_83(n7_adj_3952), .n7_adj_84(n7_adj_3951), 
            .n7_adj_85(n7_adj_3950), .n7_adj_86(n7_adj_3949), .n7_adj_87(n7_adj_3948), 
            .n7_adj_88(n7_adj_3947), .n7_adj_89(n7_adj_3946), .n7_adj_90(n7_adj_3945), 
            .n7_adj_91(n7_adj_3944), .n7_adj_92(n7_adj_3943), .n7_adj_93(n7_adj_3942), 
            .n7_adj_94(n7_adj_3941), .LM32DEBUG_ACK_O(LM32DEBUG_ACK_O), 
            .w_result({w_result}), .w_clk_cpu(w_clk_cpu), .data_bus_error_exception_N_1225(data_bus_error_exception_N_1225), 
            .n42726(n42726), .read_idx_0_d({read_idx_0_d}), .n23059(n23059), 
            .n23091(n23091), .n23058(n23058), .n23090(n23090), .n23067(n23067), 
            .n23099(n23099), .LM32D_CYC_O(LM32D_CYC_O), .n23068(n23068), 
            .n23100(n23100), .LM32I_CYC_O(LM32I_CYC_O), .n42734(n42734), 
            .n42738(n42738), .read_idx_1_d({read_idx_1_d}), .n23069(n23069), 
            .n23101(n23101), .n42732(n42732), .n23070(n23070), .n23102(n23102), 
            .n23071(n23071), .n23103(n23103), .n23072(n23072), .n23104(n23104), 
            .\counter[2] (\counter[2]_adj_101 ), .n41470(n41470), .write_idx_w({write_idx_w}), 
            .n23185(n23185), .n23186(n23186), .n23073(n23073), .n23105(n23105), 
            .n23074(n23074), .n23106(n23106), .n23075(n23075), .n23107(n23107), 
            .n23076(n23076), .n23108(n23108), .n22885(n22885), .wb_load_complete_N_2129(wb_load_complete_N_2129), 
            .reg_data_1({reg_data_1}), .n23056(n23056), .n23088(n23088), 
            .n23057(n23057), .n23089(n23089), .n22999(n22999), .n22877(n22877), 
            .n22874(n22874), .n23053(n23053), .n23085(n23085), .n23054(n23054), 
            .n23086(n23086), .n23060(n23060), .n23092(n23092), .n23061(n23061), 
            .n23093(n23093), .n23062(n23062), .n23094(n23094), .n23063(n23063), 
            .n23095(n23095), .n23064(n23064), .n23096(n23096), .n23065(n23065), 
            .n23097(n23097), .n23066(n23066), .n23098(n23098), .n23052(n23052), 
            .n23084(n23084), .n23055(n23055), .n23087(n23087), .n23077(n23077), 
            .n23109(n23109), .n23078(n23078), .n23110(n23110), .n23079(n23079), 
            .n23111(n23111), .n23080(n23080), .n23112(n23112), .n23081(n23081), 
            .n23113(n23113), .n23082(n23082), .n23114(n23114), .n23083(n23083), 
            .n23115(n23115), .i_cyc_o_N_1759(i_cyc_o_N_1759), .LM32D_WE_O(LM32D_WE_O), 
            .LM32D_DAT_O({LM32D_DAT_O}), .SHAREDBUS_DAT_O({SHAREDBUS_DAT_O}), 
            .LM32D_ADR_O({LM32D_ADR_O}), .LM32D_SEL_O({LM32D_SEL_O}), .LM32D_STB_O(LM32D_STB_O), 
            .\LM32I_ADR_O[2] (LM32I_ADR_O[2]), .\selected_1__N_344[0] (selected_1__N_344[0]), 
            .\LM32I_ADR_O[31] (LM32I_ADR_O[31]), .bus_error_f_N_1764(bus_error_f_N_1764), 
            .\LM32I_ADR_O[30] (LM32I_ADR_O[30]), .\LM32I_ADR_O[29] (LM32I_ADR_O[29]), 
            .\LM32I_ADR_O[28] (LM32I_ADR_O[28]), .\LM32I_ADR_O[27] (LM32I_ADR_O[27]), 
            .\LM32I_ADR_O[26] (LM32I_ADR_O[26]), .\LM32I_ADR_O[25] (LM32I_ADR_O[25]), 
            .\LM32I_ADR_O[24] (LM32I_ADR_O[24]), .\LM32I_ADR_O[23] (LM32I_ADR_O[23]), 
            .\LM32I_ADR_O[22] (LM32I_ADR_O[22]), .\LM32I_ADR_O[21] (LM32I_ADR_O[21]), 
            .\LM32I_ADR_O[20] (LM32I_ADR_O[20]), .\LM32I_ADR_O[19] (LM32I_ADR_O[19]), 
            .\LM32I_ADR_O[18] (LM32I_ADR_O[18]), .\LM32I_ADR_O[17] (LM32I_ADR_O[17]), 
            .\LM32I_ADR_O[16] (LM32I_ADR_O[16]), .\LM32I_ADR_O[15] (LM32I_ADR_O[15]), 
            .\LM32I_ADR_O[14] (LM32I_ADR_O[14]), .\LM32I_ADR_O[13] (LM32I_ADR_O[13]), 
            .\LM32I_ADR_O[12] (LM32I_ADR_O[12]), .\LM32I_ADR_O[11] (LM32I_ADR_O[11]), 
            .\LM32I_ADR_O[10] (LM32I_ADR_O[10]), .\LM32I_ADR_O[9] (LM32I_ADR_O[9]), 
            .\LM32I_ADR_O[8] (LM32I_ADR_O[8]), .\LM32I_ADR_O[7] (LM32I_ADR_O[7]), 
            .\LM32I_ADR_O[6] (LM32I_ADR_O[6]), .\LM32I_ADR_O[5] (LM32I_ADR_O[5]), 
            .\LM32I_ADR_O[4] (LM32I_ADR_O[4]), .\LM32I_ADR_O[3] (LM32I_ADR_O[3]), 
            .n41479(n41479), .n38871(n38871), .\data[31] (data[31]), .n87({n87}), 
            .\SHAREDBUS_SEL_I[1] (SHAREDBUS_SEL_I[1]), .n41490(n41490), 
            .\data[21] (data[21]), .\data[19] (data[19]), .w_clk_cpu_enable_303(w_clk_cpu_enable_303), 
            .\data[30] (data[30]), .n41426(n41426), .\data[29] (data[29]), 
            .\data[28] (data[28]), .n93({n4}), .n92({n1}), .n41422(n41422), 
            .n35(n35), .\data[27] (data[27]), .\data[26] (data[26]), .\data[25] (data[25]), 
            .\data[18] (data[18]), .\data[24] (data[24]), .\data[23] (data[23]), 
            .\data[17] (data[17]), .\data[16] (data[16]), .n96({n96}), 
            .\data[22] (data[22]), .\data[20] (data[20]), .\SHAREDBUS_ADR_I[10] (SHAREDBUS_ADR_I[10]), 
            .\SHAREDBUS_ADR_I[9] (SHAREDBUS_ADR_I[9]), .\SHAREDBUS_ADR_I[8] (SHAREDBUS_ADR_I[8]), 
            .\SHAREDBUS_ADR_I[7] (SHAREDBUS_ADR_I[7]), .\SHAREDBUS_ADR_I[6] (SHAREDBUS_ADR_I[6]), 
            .\SHAREDBUS_ADR_I[5] (SHAREDBUS_ADR_I[5]), .\SHAREDBUS_ADR_I[4] (SHAREDBUS_ADR_I[4]), 
            .\SHAREDBUS_ADR_I[3] (SHAREDBUS_ADR_I[3]), .\SHAREDBUS_ADR_I[2] (SHAREDBUS_ADR_I[2]), 
            .VCC_net(VCC_net), .counter_2__N_178(counter_2__N_178)) /* synthesis syn_module_defined=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(519[2] 560[36])
    
endmodule
//
// Verilog Description of module \asram_top(SRAM_DATA_WIDTH=8,SRAM_ADDR_WIDTH=19,SRAM_BE_WIDTH=1,READ_LATENCY=2,WRITE_LATENCY=2,DATA_OUTPUT_REG=1) 
//

module \asram_top(SRAM_DATA_WIDTH=8,SRAM_ADDR_WIDTH=19,SRAM_BE_WIDTH=1,READ_LATENCY=2,WRITE_LATENCY=2,DATA_OUTPUT_REG=1)  (sramASRAM_DAT_O, 
            sramsram_data_in, n21531, n41405, n7, n41393, n36822, 
            n41501, n7_adj_100, n41356, \SHAREDBUS_SEL_I[1] , n41344, 
            w_clk_cpu, tmp_ack_o, n41488, n24342, n28684, sram_adr_c_0, 
            \genblk5.tmp_ack_o_d , n42723, sramsram_data_out, w_clk_cpu_enable_900, 
            n26128, sram_adr_c_18, \SHAREDBUS_ADR_I[18] , sram_adr_c_17, 
            \SHAREDBUS_ADR_I[17] , sram_adr_c_16, \SHAREDBUS_ADR_I[16] , 
            sram_adr_c_15, \SHAREDBUS_ADR_I[15] , \SHAREDBUS_ADR_I[0] , 
            sram_adr_c_14, \SHAREDBUS_ADR_I[14] , sram_adr_c_13, n41435, 
            \LM32D_ADR_O[1] , n41412, sram_adr_c_12, \SHAREDBUS_ADR_I[12] , 
            sram_adr_c_11, \SHAREDBUS_ADR_I[11] , sram_adr_c_10, \SHAREDBUS_ADR_I[10] , 
            sram_adr_c_9, \SHAREDBUS_ADR_I[9] , n41353, sram_adr_c_8, 
            \SHAREDBUS_ADR_I[8] , sram_adr_c_7, \SHAREDBUS_ADR_I[7] , 
            sram_adr_c_6, \SHAREDBUS_ADR_I[6] , sram_adr_c_5, \SHAREDBUS_ADR_I[5] , 
            sram_adr_c_4, \SHAREDBUS_ADR_I[4] , sram_adr_c_3, \SHAREDBUS_ADR_I[3] , 
            sram_adr_c_2, \SHAREDBUS_ADR_I[2] , sram_adr_c_1, LM32D_SEL_O, 
            selected, n41424, n38761, PIO_OUT_7__N_3327, n41423, n41490, 
            n25515, n25664, w_clk_cpu_enable_303, n41363, n24709, 
            n39016, LM32D_DAT_O, n36688, n183, n22230, n38998, n31536, 
            sram_data_out_nxt_7__N_3203, n37005, n39018, n40734, state_nxt_1__N_3154, 
            n41429, n41390, n40733, n41453, n41392, n41479, n41469, 
            n41455, \data[28] , \SHAREDBUS_DAT_I[28] , n96, \data[29] , 
            \SHAREDBUS_DAT_I[29] , \data[30] , \SHAREDBUS_DAT_I[30] , 
            \data[31] , \SHAREDBUS_DAT_I[31] , \data[27] , \SHAREDBUS_DAT_I[27] , 
            \data[26] , \SHAREDBUS_DAT_I[26] , \data[25] , \SHAREDBUS_DAT_I[25] , 
            \data[24] , \SHAREDBUS_DAT_I[24] , \tmp_dat_o_nxt_31__N_3207[19] , 
            LM32D_WE_O, sram_oen_c, n41426) /* synthesis syn_module_defined=1 */ ;
    output [31:0]sramASRAM_DAT_O;
    input [7:0]sramsram_data_in;
    output n21531;
    input n41405;
    output n7;
    input n41393;
    input n36822;
    output n41501;
    output n7_adj_100;
    input n41356;
    input \SHAREDBUS_SEL_I[1] ;
    output n41344;
    input w_clk_cpu;
    output tmp_ack_o;
    output n41488;
    input n24342;
    output n28684;
    output sram_adr_c_0;
    output \genblk5.tmp_ack_o_d ;
    output n42723;
    output [7:0]sramsram_data_out;
    output w_clk_cpu_enable_900;
    input n26128;
    output sram_adr_c_18;
    input \SHAREDBUS_ADR_I[18] ;
    output sram_adr_c_17;
    input \SHAREDBUS_ADR_I[17] ;
    output sram_adr_c_16;
    input \SHAREDBUS_ADR_I[16] ;
    output sram_adr_c_15;
    input \SHAREDBUS_ADR_I[15] ;
    input \SHAREDBUS_ADR_I[0] ;
    output sram_adr_c_14;
    input \SHAREDBUS_ADR_I[14] ;
    output sram_adr_c_13;
    input n41435;
    input \LM32D_ADR_O[1] ;
    input n41412;
    output sram_adr_c_12;
    input \SHAREDBUS_ADR_I[12] ;
    output sram_adr_c_11;
    input \SHAREDBUS_ADR_I[11] ;
    output sram_adr_c_10;
    input \SHAREDBUS_ADR_I[10] ;
    output sram_adr_c_9;
    input \SHAREDBUS_ADR_I[9] ;
    input n41353;
    output sram_adr_c_8;
    input \SHAREDBUS_ADR_I[8] ;
    output sram_adr_c_7;
    input \SHAREDBUS_ADR_I[7] ;
    output sram_adr_c_6;
    input \SHAREDBUS_ADR_I[6] ;
    output sram_adr_c_5;
    input \SHAREDBUS_ADR_I[5] ;
    output sram_adr_c_4;
    input \SHAREDBUS_ADR_I[4] ;
    output sram_adr_c_3;
    input \SHAREDBUS_ADR_I[3] ;
    output sram_adr_c_2;
    input \SHAREDBUS_ADR_I[2] ;
    output sram_adr_c_1;
    input [3:0]LM32D_SEL_O;
    input [1:0]selected;
    output n41424;
    input n38761;
    output PIO_OUT_7__N_3327;
    input n41423;
    input n41490;
    output n25515;
    output n25664;
    input w_clk_cpu_enable_303;
    input n41363;
    output n24709;
    output n39016;
    input [31:0]LM32D_DAT_O;
    input n36688;
    input n183;
    input n22230;
    input n38998;
    input n31536;
    input sram_data_out_nxt_7__N_3203;
    input n37005;
    input n39018;
    input n40734;
    input state_nxt_1__N_3154;
    input n41429;
    input n41390;
    output n40733;
    output n41453;
    input n41392;
    input n41479;
    input n41469;
    input n41455;
    input \data[28] ;
    input \SHAREDBUS_DAT_I[28] ;
    output [7:0]n96;
    input \data[29] ;
    input \SHAREDBUS_DAT_I[29] ;
    input \data[30] ;
    input \SHAREDBUS_DAT_I[30] ;
    input \data[31] ;
    input \SHAREDBUS_DAT_I[31] ;
    input \data[27] ;
    input \SHAREDBUS_DAT_I[27] ;
    input \data[26] ;
    input \SHAREDBUS_DAT_I[26] ;
    input \data[25] ;
    input \SHAREDBUS_DAT_I[25] ;
    input \data[24] ;
    input \SHAREDBUS_DAT_I[24] ;
    input \tmp_dat_o_nxt_31__N_3207[19] ;
    input LM32D_WE_O;
    output sram_oen_c;
    input n41426;
    
    wire w_clk_cpu /* synthesis SET_AS_NETWORK=w_clk_cpu, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(22[6:15])
    
    \asram_core(SRAM_DATA_WIDTH=8,SRAM_ADDR_WIDTH=19,SRAM_BE_WIDTH=1,READ_LATENCY=2,WRITE_LATENCY=2,DATA_OUTPUT_REG=1)  core_inst (.sramASRAM_DAT_O({sramASRAM_DAT_O}), 
            .sramsram_data_in({sramsram_data_in}), .n21531(n21531), .n41405(n41405), 
            .n7(n7), .n41393(n41393), .n36822(n36822), .n41501(n41501), 
            .n7_adj_99(n7_adj_100), .n41356(n41356), .\SHAREDBUS_SEL_I[1] (\SHAREDBUS_SEL_I[1] ), 
            .n41344(n41344), .w_clk_cpu(w_clk_cpu), .tmp_ack_o(tmp_ack_o), 
            .n41488(n41488), .n24342(n24342), .n28684(n28684), .sram_adr_c_0(sram_adr_c_0), 
            .\genblk5.tmp_ack_o_d (\genblk5.tmp_ack_o_d ), .n42723(n42723), 
            .sramsram_data_out({sramsram_data_out}), .w_clk_cpu_enable_900(w_clk_cpu_enable_900), 
            .n26128(n26128), .sram_adr_c_18(sram_adr_c_18), .\SHAREDBUS_ADR_I[18] (\SHAREDBUS_ADR_I[18] ), 
            .sram_adr_c_17(sram_adr_c_17), .\SHAREDBUS_ADR_I[17] (\SHAREDBUS_ADR_I[17] ), 
            .sram_adr_c_16(sram_adr_c_16), .\SHAREDBUS_ADR_I[16] (\SHAREDBUS_ADR_I[16] ), 
            .sram_adr_c_15(sram_adr_c_15), .\SHAREDBUS_ADR_I[15] (\SHAREDBUS_ADR_I[15] ), 
            .\SHAREDBUS_ADR_I[0] (\SHAREDBUS_ADR_I[0] ), .sram_adr_c_14(sram_adr_c_14), 
            .\SHAREDBUS_ADR_I[14] (\SHAREDBUS_ADR_I[14] ), .sram_adr_c_13(sram_adr_c_13), 
            .n41435(n41435), .\LM32D_ADR_O[1] (\LM32D_ADR_O[1] ), .n41412(n41412), 
            .sram_adr_c_12(sram_adr_c_12), .\SHAREDBUS_ADR_I[12] (\SHAREDBUS_ADR_I[12] ), 
            .sram_adr_c_11(sram_adr_c_11), .\SHAREDBUS_ADR_I[11] (\SHAREDBUS_ADR_I[11] ), 
            .sram_adr_c_10(sram_adr_c_10), .\SHAREDBUS_ADR_I[10] (\SHAREDBUS_ADR_I[10] ), 
            .sram_adr_c_9(sram_adr_c_9), .\SHAREDBUS_ADR_I[9] (\SHAREDBUS_ADR_I[9] ), 
            .n41353(n41353), .sram_adr_c_8(sram_adr_c_8), .\SHAREDBUS_ADR_I[8] (\SHAREDBUS_ADR_I[8] ), 
            .sram_adr_c_7(sram_adr_c_7), .\SHAREDBUS_ADR_I[7] (\SHAREDBUS_ADR_I[7] ), 
            .sram_adr_c_6(sram_adr_c_6), .\SHAREDBUS_ADR_I[6] (\SHAREDBUS_ADR_I[6] ), 
            .sram_adr_c_5(sram_adr_c_5), .\SHAREDBUS_ADR_I[5] (\SHAREDBUS_ADR_I[5] ), 
            .sram_adr_c_4(sram_adr_c_4), .\SHAREDBUS_ADR_I[4] (\SHAREDBUS_ADR_I[4] ), 
            .sram_adr_c_3(sram_adr_c_3), .\SHAREDBUS_ADR_I[3] (\SHAREDBUS_ADR_I[3] ), 
            .sram_adr_c_2(sram_adr_c_2), .\SHAREDBUS_ADR_I[2] (\SHAREDBUS_ADR_I[2] ), 
            .sram_adr_c_1(sram_adr_c_1), .LM32D_SEL_O({LM32D_SEL_O}), .selected({selected}), 
            .n41424(n41424), .n38761(n38761), .PIO_OUT_7__N_3327(PIO_OUT_7__N_3327), 
            .n41423(n41423), .n41490(n41490), .n25515(n25515), .n25664(n25664), 
            .w_clk_cpu_enable_303(w_clk_cpu_enable_303), .n41363(n41363), 
            .n24709(n24709), .n39016(n39016), .LM32D_DAT_O({LM32D_DAT_O}), 
            .n36688(n36688), .n183(n183), .n22230(n22230), .n38998(n38998), 
            .n31536(n31536), .sram_data_out_nxt_7__N_3203(sram_data_out_nxt_7__N_3203), 
            .n37005(n37005), .n39018(n39018), .n40734(n40734), .state_nxt_1__N_3154(state_nxt_1__N_3154), 
            .n41429(n41429), .n41390(n41390), .n40733(n40733), .n41453(n41453), 
            .n41392(n41392), .n41479(n41479), .n41469(n41469), .n41455(n41455), 
            .\data[28] (\data[28] ), .\SHAREDBUS_DAT_I[28] (\SHAREDBUS_DAT_I[28] ), 
            .n96({n96}), .\data[29] (\data[29] ), .\SHAREDBUS_DAT_I[29] (\SHAREDBUS_DAT_I[29] ), 
            .\data[30] (\data[30] ), .\SHAREDBUS_DAT_I[30] (\SHAREDBUS_DAT_I[30] ), 
            .\data[31] (\data[31] ), .\SHAREDBUS_DAT_I[31] (\SHAREDBUS_DAT_I[31] ), 
            .\data[27] (\data[27] ), .\SHAREDBUS_DAT_I[27] (\SHAREDBUS_DAT_I[27] ), 
            .\data[26] (\data[26] ), .\SHAREDBUS_DAT_I[26] (\SHAREDBUS_DAT_I[26] ), 
            .\data[25] (\data[25] ), .\SHAREDBUS_DAT_I[25] (\SHAREDBUS_DAT_I[25] ), 
            .\data[24] (\data[24] ), .\SHAREDBUS_DAT_I[24] (\SHAREDBUS_DAT_I[24] ), 
            .\tmp_dat_o_nxt_31__N_3207[19] (\tmp_dat_o_nxt_31__N_3207[19] ), 
            .LM32D_WE_O(LM32D_WE_O), .sram_oen_c(sram_oen_c), .n41426(n41426)) /* synthesis syn_module_defined=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_top.v(109[4] 128[36])
    
endmodule
//
// Verilog Description of module \asram_core(SRAM_DATA_WIDTH=8,SRAM_ADDR_WIDTH=19,SRAM_BE_WIDTH=1,READ_LATENCY=2,WRITE_LATENCY=2,DATA_OUTPUT_REG=1) 
//

module \asram_core(SRAM_DATA_WIDTH=8,SRAM_ADDR_WIDTH=19,SRAM_BE_WIDTH=1,READ_LATENCY=2,WRITE_LATENCY=2,DATA_OUTPUT_REG=1)  (sramASRAM_DAT_O, 
            sramsram_data_in, n21531, n41405, n7, n41393, n36822, 
            n41501, n7_adj_99, n41356, \SHAREDBUS_SEL_I[1] , n41344, 
            w_clk_cpu, tmp_ack_o, n41488, n24342, n28684, sram_adr_c_0, 
            \genblk5.tmp_ack_o_d , n42723, sramsram_data_out, w_clk_cpu_enable_900, 
            n26128, sram_adr_c_18, \SHAREDBUS_ADR_I[18] , sram_adr_c_17, 
            \SHAREDBUS_ADR_I[17] , sram_adr_c_16, \SHAREDBUS_ADR_I[16] , 
            sram_adr_c_15, \SHAREDBUS_ADR_I[15] , \SHAREDBUS_ADR_I[0] , 
            sram_adr_c_14, \SHAREDBUS_ADR_I[14] , sram_adr_c_13, n41435, 
            \LM32D_ADR_O[1] , n41412, sram_adr_c_12, \SHAREDBUS_ADR_I[12] , 
            sram_adr_c_11, \SHAREDBUS_ADR_I[11] , sram_adr_c_10, \SHAREDBUS_ADR_I[10] , 
            sram_adr_c_9, \SHAREDBUS_ADR_I[9] , n41353, sram_adr_c_8, 
            \SHAREDBUS_ADR_I[8] , sram_adr_c_7, \SHAREDBUS_ADR_I[7] , 
            sram_adr_c_6, \SHAREDBUS_ADR_I[6] , sram_adr_c_5, \SHAREDBUS_ADR_I[5] , 
            sram_adr_c_4, \SHAREDBUS_ADR_I[4] , sram_adr_c_3, \SHAREDBUS_ADR_I[3] , 
            sram_adr_c_2, \SHAREDBUS_ADR_I[2] , sram_adr_c_1, LM32D_SEL_O, 
            selected, n41424, n38761, PIO_OUT_7__N_3327, n41423, n41490, 
            n25515, n25664, w_clk_cpu_enable_303, n41363, n24709, 
            n39016, LM32D_DAT_O, n36688, n183, n22230, n38998, n31536, 
            sram_data_out_nxt_7__N_3203, n37005, n39018, n40734, state_nxt_1__N_3154, 
            n41429, n41390, n40733, n41453, n41392, n41479, n41469, 
            n41455, \data[28] , \SHAREDBUS_DAT_I[28] , n96, \data[29] , 
            \SHAREDBUS_DAT_I[29] , \data[30] , \SHAREDBUS_DAT_I[30] , 
            \data[31] , \SHAREDBUS_DAT_I[31] , \data[27] , \SHAREDBUS_DAT_I[27] , 
            \data[26] , \SHAREDBUS_DAT_I[26] , \data[25] , \SHAREDBUS_DAT_I[25] , 
            \data[24] , \SHAREDBUS_DAT_I[24] , \tmp_dat_o_nxt_31__N_3207[19] , 
            LM32D_WE_O, sram_oen_c, n41426) /* synthesis syn_module_defined=1 */ ;
    output [31:0]sramASRAM_DAT_O;
    input [7:0]sramsram_data_in;
    output n21531;
    input n41405;
    output n7;
    input n41393;
    input n36822;
    output n41501;
    output n7_adj_99;
    input n41356;
    input \SHAREDBUS_SEL_I[1] ;
    output n41344;
    input w_clk_cpu;
    output tmp_ack_o;
    output n41488;
    input n24342;
    output n28684;
    output sram_adr_c_0;
    output \genblk5.tmp_ack_o_d ;
    output n42723;
    output [7:0]sramsram_data_out;
    output w_clk_cpu_enable_900;
    input n26128;
    output sram_adr_c_18;
    input \SHAREDBUS_ADR_I[18] ;
    output sram_adr_c_17;
    input \SHAREDBUS_ADR_I[17] ;
    output sram_adr_c_16;
    input \SHAREDBUS_ADR_I[16] ;
    output sram_adr_c_15;
    input \SHAREDBUS_ADR_I[15] ;
    input \SHAREDBUS_ADR_I[0] ;
    output sram_adr_c_14;
    input \SHAREDBUS_ADR_I[14] ;
    output sram_adr_c_13;
    input n41435;
    input \LM32D_ADR_O[1] ;
    input n41412;
    output sram_adr_c_12;
    input \SHAREDBUS_ADR_I[12] ;
    output sram_adr_c_11;
    input \SHAREDBUS_ADR_I[11] ;
    output sram_adr_c_10;
    input \SHAREDBUS_ADR_I[10] ;
    output sram_adr_c_9;
    input \SHAREDBUS_ADR_I[9] ;
    input n41353;
    output sram_adr_c_8;
    input \SHAREDBUS_ADR_I[8] ;
    output sram_adr_c_7;
    input \SHAREDBUS_ADR_I[7] ;
    output sram_adr_c_6;
    input \SHAREDBUS_ADR_I[6] ;
    output sram_adr_c_5;
    input \SHAREDBUS_ADR_I[5] ;
    output sram_adr_c_4;
    input \SHAREDBUS_ADR_I[4] ;
    output sram_adr_c_3;
    input \SHAREDBUS_ADR_I[3] ;
    output sram_adr_c_2;
    input \SHAREDBUS_ADR_I[2] ;
    output sram_adr_c_1;
    input [3:0]LM32D_SEL_O;
    input [1:0]selected;
    output n41424;
    input n38761;
    output PIO_OUT_7__N_3327;
    input n41423;
    input n41490;
    output n25515;
    output n25664;
    input w_clk_cpu_enable_303;
    input n41363;
    output n24709;
    output n39016;
    input [31:0]LM32D_DAT_O;
    input n36688;
    input n183;
    input n22230;
    input n38998;
    input n31536;
    input sram_data_out_nxt_7__N_3203;
    input n37005;
    input n39018;
    input n40734;
    input state_nxt_1__N_3154;
    input n41429;
    input n41390;
    output n40733;
    output n41453;
    input n41392;
    input n41479;
    input n41469;
    input n41455;
    input \data[28] ;
    input \SHAREDBUS_DAT_I[28] ;
    output [7:0]n96;
    input \data[29] ;
    input \SHAREDBUS_DAT_I[29] ;
    input \data[30] ;
    input \SHAREDBUS_DAT_I[30] ;
    input \data[31] ;
    input \SHAREDBUS_DAT_I[31] ;
    input \data[27] ;
    input \SHAREDBUS_DAT_I[27] ;
    input \data[26] ;
    input \SHAREDBUS_DAT_I[26] ;
    input \data[25] ;
    input \SHAREDBUS_DAT_I[25] ;
    input \data[24] ;
    input \SHAREDBUS_DAT_I[24] ;
    input \tmp_dat_o_nxt_31__N_3207[19] ;
    input LM32D_WE_O;
    output sram_oen_c;
    input n41426;
    
    wire w_clk_cpu /* synthesis SET_AS_NETWORK=w_clk_cpu, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(22[6:15])
    wire [1:0]cycle;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(101[16:21])
    wire [15:0]n21518;
    wire [31:0]n467;
    wire [31:0]tmp_dat_o_nxt_31__N_3094;
    
    wire cycle_counter_nxt_1__N_3179, w_clk_cpu_enable_349, n41343, n41342;
    wire [1:0]state;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(111[14:19])
    
    wire n5, n23818, tmp_ack_o_nxt_N_3277, w_clk_cpu_enable_648;
    wire [3:0]dly;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(108[21:24])
    
    wire n633;
    wire [3:0]dly_nxt_3__N_3165;
    wire [31:0]tmp_dat_o_nxt_31__N_3207;
    wire [1:0]cycle_counter_nxt;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(109[44:61])
    
    wire w_clk_cpu_enable_339;
    wire [18:0]sram_addr_nxt;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(103[30:43])
    
    wire w_clk_cpu_enable_184, n1, n39070, n26089, n26105, n39339, 
        n26111, n26073, n26087, n26103, n26071, n26085, n26101, 
        n26069, n26083, n26099, n26093, n26109, n26115, n26091, 
        n26107, n26113, n26067, n26081, n26097, n26045, n26047, 
        n26049, sram_addr_nxt_18__N_3187, sram_addr_nxt_18__N_3069, n41478, 
        n26018;
    wire [1:0]cycle_counter_nxt_1__N_3177;
    wire [1:0]acycle;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(109[21:27])
    
    wire tmp_dat_o_nxt_31__N_3127, n29457, n29460, w_clk_cpu_enable_363;
    wire [3:0]dly_nxt;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(108[26:33])
    
    wire dly_nxt_3__N_3169, n41500, sram_data_out_nxt_7__N_3086, n41497, 
        sram_data_out_nxt_7__N_3201, n41374, n5_adj_3938, n41496, n14;
    wire [31:0]tmp_dat_o_nxt_31__N_3239;
    
    wire w_clk_cpu_enable_527, n38992, w_clk_cpu_enable_566, n41618, 
        w_clk_cpu_enable_577, w_clk_cpu_enable_619, n41341, n41445, 
        n41619, n36806;
    
    LUT4 mux_19179_i6_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(sramASRAM_DAT_O[21]), 
         .D(sramsram_data_in[5]), .Z(n21518[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam mux_19179_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19179_i4_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(sramASRAM_DAT_O[19]), 
         .D(sramsram_data_in[3]), .Z(n21531)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam mux_19179_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19179_i3_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(sramASRAM_DAT_O[18]), 
         .D(sramsram_data_in[2]), .Z(n21518[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam mux_19179_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19179_i2_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(sramASRAM_DAT_O[17]), 
         .D(sramsram_data_in[1]), .Z(n21518[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam mux_19179_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 tmp_dat_o_nxt_31__I_151_i15_4_lut (.A(sramsram_data_in[6]), .B(n467[14]), 
         .C(n41405), .D(n7), .Z(tmp_dat_o_nxt_31__N_3094[14])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i15_4_lut.init = 16'hca0a;
    LUT4 mux_199_i15_4_lut (.A(n21518[14]), .B(sramsram_data_in[6]), .C(n41393), 
         .D(n36822), .Z(n467[14])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(555[10] 562[17])
    defparam mux_199_i15_4_lut.init = 16'h0aca;
    LUT4 tmp_dat_o_nxt_31__I_151_i14_4_lut (.A(sramsram_data_in[5]), .B(n467[13]), 
         .C(n41405), .D(n7), .Z(tmp_dat_o_nxt_31__N_3094[13])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i14_4_lut.init = 16'hca0a;
    LUT4 mux_199_i14_4_lut (.A(n21518[13]), .B(sramsram_data_in[5]), .C(n41393), 
         .D(n36822), .Z(n467[13])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(555[10] 562[17])
    defparam mux_199_i14_4_lut.init = 16'h0aca;
    LUT4 i1_2_lut_4_lut (.A(n41501), .B(n7_adj_99), .C(n41356), .D(cycle_counter_nxt_1__N_3179), 
         .Z(w_clk_cpu_enable_349)) /* synthesis lut_function=((B (D)+!B (C+(D)))+!A) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(204[9:95])
    defparam i1_2_lut_4_lut.init = 16'hff75;
    LUT4 tmp_dat_o_nxt_31__I_151_i13_4_lut (.A(sramsram_data_in[4]), .B(n467[12]), 
         .C(n41405), .D(n7), .Z(tmp_dat_o_nxt_31__N_3094[12])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i13_4_lut.init = 16'hca0a;
    LUT4 mux_199_i13_4_lut (.A(n21518[12]), .B(sramsram_data_in[4]), .C(n41393), 
         .D(n36822), .Z(n467[12])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(555[10] 562[17])
    defparam mux_199_i13_4_lut.init = 16'h0aca;
    LUT4 tmp_dat_o_nxt_31__I_151_i12_4_lut (.A(sramsram_data_in[3]), .B(n467[11]), 
         .C(n41405), .D(n7), .Z(tmp_dat_o_nxt_31__N_3094[11])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i12_4_lut.init = 16'hca0a;
    PFUMX i38565 (.BLUT(n41343), .ALUT(n41342), .C0(\SHAREDBUS_SEL_I[1] ), 
          .Z(n41344));
    LUT4 mux_199_i12_4_lut (.A(n21518[11]), .B(sramsram_data_in[3]), .C(n41393), 
         .D(n36822), .Z(n467[11])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(555[10] 562[17])
    defparam mux_199_i12_4_lut.init = 16'h0aca;
    FD1S3IX state_i1 (.D(n23818), .CK(w_clk_cpu), .CD(n5), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam state_i1.GSR = "ENABLED";
    LUT4 tmp_dat_o_nxt_31__I_151_i11_4_lut (.A(sramsram_data_in[2]), .B(n467[10]), 
         .C(n41405), .D(n7), .Z(tmp_dat_o_nxt_31__N_3094[10])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i11_4_lut.init = 16'hca0a;
    LUT4 mux_199_i11_4_lut (.A(n21518[10]), .B(sramsram_data_in[2]), .C(n41393), 
         .D(n36822), .Z(n467[10])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(555[10] 562[17])
    defparam mux_199_i11_4_lut.init = 16'h0aca;
    FD1S3IX tmp_ack_o_248 (.D(tmp_ack_o_nxt_N_3277), .CK(w_clk_cpu), .CD(n41488), 
            .Q(tmp_ack_o));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(669[4:34])
    defparam tmp_ack_o_248.GSR = "ENABLED";
    LUT4 tmp_dat_o_nxt_31__I_151_i10_4_lut (.A(sramsram_data_in[1]), .B(n467[9]), 
         .C(n41405), .D(n7), .Z(tmp_dat_o_nxt_31__N_3094[9])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i10_4_lut.init = 16'hca0a;
    LUT4 mux_199_i10_4_lut (.A(n21518[9]), .B(sramsram_data_in[1]), .C(n41393), 
         .D(n36822), .Z(n467[9])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(555[10] 562[17])
    defparam mux_199_i10_4_lut.init = 16'h0aca;
    LUT4 tmp_dat_o_nxt_31__I_151_i9_4_lut (.A(sramsram_data_in[0]), .B(n467[8]), 
         .C(n41405), .D(n7), .Z(tmp_dat_o_nxt_31__N_3094[8])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i9_4_lut.init = 16'hca0a;
    LUT4 mux_199_i9_4_lut (.A(n21518[8]), .B(sramsram_data_in[0]), .C(n41393), 
         .D(n36822), .Z(n467[8])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(555[10] 562[17])
    defparam mux_199_i9_4_lut.init = 16'h0aca;
    LUT4 tmp_dat_o_nxt_31__I_151_i8_4_lut (.A(sramsram_data_in[7]), .B(n467[7]), 
         .C(n41405), .D(n7), .Z(tmp_dat_o_nxt_31__N_3094[7])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i8_4_lut.init = 16'hca0a;
    LUT4 mux_199_i8_4_lut (.A(n21518[7]), .B(sramsram_data_in[7]), .C(n41393), 
         .D(n24342), .Z(n467[7])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(555[10] 562[17])
    defparam mux_199_i8_4_lut.init = 16'hca0a;
    LUT4 tmp_dat_o_nxt_31__I_151_i7_4_lut (.A(sramsram_data_in[6]), .B(n467[6]), 
         .C(n41405), .D(n7), .Z(tmp_dat_o_nxt_31__N_3094[6])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i7_4_lut.init = 16'hca0a;
    LUT4 mux_199_i7_4_lut (.A(n21518[6]), .B(sramsram_data_in[6]), .C(n41393), 
         .D(n24342), .Z(n467[6])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(555[10] 562[17])
    defparam mux_199_i7_4_lut.init = 16'hca0a;
    LUT4 tmp_dat_o_nxt_31__I_151_i6_4_lut (.A(sramsram_data_in[5]), .B(n467[5]), 
         .C(n41405), .D(n7), .Z(tmp_dat_o_nxt_31__N_3094[5])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i6_4_lut.init = 16'hca0a;
    LUT4 mux_199_i6_4_lut (.A(n21518[5]), .B(sramsram_data_in[5]), .C(n41393), 
         .D(n24342), .Z(n467[5])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(555[10] 562[17])
    defparam mux_199_i6_4_lut.init = 16'hca0a;
    LUT4 tmp_dat_o_nxt_31__I_151_i5_4_lut (.A(sramsram_data_in[4]), .B(n467[4]), 
         .C(n41405), .D(n7), .Z(tmp_dat_o_nxt_31__N_3094[4])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i5_4_lut.init = 16'hca0a;
    LUT4 mux_199_i5_4_lut (.A(n21518[4]), .B(sramsram_data_in[4]), .C(n41393), 
         .D(n24342), .Z(n467[4])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(555[10] 562[17])
    defparam mux_199_i5_4_lut.init = 16'hca0a;
    LUT4 tmp_dat_o_nxt_31__I_151_i4_4_lut (.A(sramsram_data_in[3]), .B(n467[3]), 
         .C(n41405), .D(n7), .Z(tmp_dat_o_nxt_31__N_3094[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i4_4_lut.init = 16'hca0a;
    LUT4 i20886_1_lut (.A(state[0]), .Z(n5)) /* synthesis lut_function=(!(A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(535[12:28])
    defparam i20886_1_lut.init = 16'h5555;
    LUT4 mux_199_i4_4_lut (.A(n21531), .B(sramsram_data_in[3]), .C(n41393), 
         .D(n24342), .Z(n467[3])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(555[10] 562[17])
    defparam mux_199_i4_4_lut.init = 16'hca0a;
    LUT4 tmp_dat_o_nxt_31__I_151_i3_4_lut (.A(sramsram_data_in[2]), .B(n467[2]), 
         .C(n41405), .D(n7), .Z(tmp_dat_o_nxt_31__N_3094[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i3_4_lut.init = 16'hca0a;
    LUT4 mux_199_i3_4_lut (.A(n21518[2]), .B(sramsram_data_in[2]), .C(n41393), 
         .D(n24342), .Z(n467[2])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(555[10] 562[17])
    defparam mux_199_i3_4_lut.init = 16'hca0a;
    LUT4 tmp_dat_o_nxt_31__I_151_i2_4_lut (.A(sramsram_data_in[1]), .B(n467[1]), 
         .C(n41405), .D(n7), .Z(tmp_dat_o_nxt_31__N_3094[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i2_4_lut.init = 16'hca0a;
    LUT4 mux_199_i2_4_lut (.A(n21518[1]), .B(sramsram_data_in[1]), .C(n41393), 
         .D(n24342), .Z(n467[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(555[10] 562[17])
    defparam mux_199_i2_4_lut.init = 16'hca0a;
    FD1P3AX tmp_dat_o_i0_i0 (.D(tmp_dat_o_nxt_31__N_3094[0]), .SP(w_clk_cpu_enable_648), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[0])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i0.GSR = "ENABLED";
    FD1S3IX dly_i0 (.D(dly_nxt_3__N_3165[0]), .CK(w_clk_cpu), .CD(n633), 
            .Q(dly[0])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam dly_i0.GSR = "ENABLED";
    LUT4 mux_200_i18_4_lut (.A(n21518[1]), .B(n28684), .C(n7), .D(sramsram_data_in[1]), 
         .Z(tmp_dat_o_nxt_31__N_3207[17])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(549[13] 562[17])
    defparam mux_200_i18_4_lut.init = 16'hca0a;
    FD1S3AX cycle_counter_i0 (.D(cycle_counter_nxt[0]), .CK(w_clk_cpu), 
            .Q(cycle[0])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(216[7:45])
    defparam cycle_counter_i0.GSR = "ENABLED";
    FD1P3AX sram_addr_i1 (.D(sram_addr_nxt[0]), .SP(w_clk_cpu_enable_339), 
            .CK(w_clk_cpu), .Q(sram_adr_c_0)) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_addr_i1.GSR = "ENABLED";
    LUT4 mux_200_i17_4_lut (.A(n21518[0]), .B(n28684), .C(n7), .D(sramsram_data_in[0]), 
         .Z(tmp_dat_o_nxt_31__N_3207[16])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(549[13] 562[17])
    defparam mux_200_i17_4_lut.init = 16'hca0a;
    FD1P3AX state_i0 (.D(n1), .SP(w_clk_cpu_enable_184), .CK(w_clk_cpu), 
            .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam state_i0.GSR = "ENABLED";
    FD1S3AX \genblk5.tmp_ack_o_d_249  (.D(tmp_ack_o), .CK(w_clk_cpu), .Q(\genblk5.tmp_ack_o_d )) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(678[7:35])
    defparam \genblk5.tmp_ack_o_d_249 .GSR = "ENABLED";
    LUT4 i3_4_lut (.A(n42723), .B(dly[0]), .C(dly[1]), .D(n39070), .Z(tmp_ack_o_nxt_N_3277)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3_4_lut.init = 16'h0010;
    PFUMX i23469 (.BLUT(n26089), .ALUT(n26105), .C0(n39339), .Z(n26111));
    LUT4 i36526_2_lut (.A(dly[2]), .B(dly[3]), .Z(n39070)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i36526_2_lut.init = 16'heeee;
    PFUMX i23461 (.BLUT(n26073), .ALUT(n26087), .C0(n39339), .Z(n26103));
    PFUMX i23459 (.BLUT(n26071), .ALUT(n26085), .C0(n39339), .Z(n26101));
    PFUMX i23457 (.BLUT(n26069), .ALUT(n26083), .C0(n39339), .Z(n26099));
    FD1P3IX sram_data_out_i1 (.D(n26103), .SP(w_clk_cpu_enable_900), .CD(n26128), 
            .CK(w_clk_cpu), .Q(sramsram_data_out[1])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_data_out_i1.GSR = "ENABLED";
    PFUMX i23473 (.BLUT(n26093), .ALUT(n26109), .C0(n39339), .Z(n26115));
    PFUMX i23471 (.BLUT(n26091), .ALUT(n26107), .C0(n39339), .Z(n26113));
    PFUMX i23455 (.BLUT(n26067), .ALUT(n26081), .C0(n39339), .Z(n26097));
    FD1P3IX sram_data_out_i2 (.D(n26101), .SP(w_clk_cpu_enable_900), .CD(n26128), 
            .CK(w_clk_cpu), .Q(sramsram_data_out[2])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_data_out_i2.GSR = "ENABLED";
    PFUMX i23408 (.BLUT(n26045), .ALUT(n26047), .C0(n39339), .Z(n26049));
    FD1P3IX sram_data_out_i3 (.D(n26099), .SP(w_clk_cpu_enable_900), .CD(n26128), 
            .CK(w_clk_cpu), .Q(sramsram_data_out[3])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_data_out_i3.GSR = "ENABLED";
    FD1P3IX sram_data_out_i4 (.D(n26097), .SP(w_clk_cpu_enable_900), .CD(n26128), 
            .CK(w_clk_cpu), .Q(sramsram_data_out[4])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_data_out_i4.GSR = "ENABLED";
    FD1P3IX sram_data_out_i5 (.D(n26115), .SP(w_clk_cpu_enable_900), .CD(n26128), 
            .CK(w_clk_cpu), .Q(sramsram_data_out[5])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_data_out_i5.GSR = "ENABLED";
    FD1P3AX sram_addr_i19 (.D(\SHAREDBUS_ADR_I[18] ), .SP(w_clk_cpu_enable_339), 
            .CK(w_clk_cpu), .Q(sram_adr_c_18)) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_addr_i19.GSR = "ENABLED";
    FD1P3AX sram_addr_i18 (.D(\SHAREDBUS_ADR_I[17] ), .SP(w_clk_cpu_enable_339), 
            .CK(w_clk_cpu), .Q(sram_adr_c_17)) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_addr_i18.GSR = "ENABLED";
    FD1P3AX sram_addr_i17 (.D(\SHAREDBUS_ADR_I[16] ), .SP(w_clk_cpu_enable_339), 
            .CK(w_clk_cpu), .Q(sram_adr_c_16)) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_addr_i17.GSR = "ENABLED";
    FD1P3AX sram_addr_i16 (.D(\SHAREDBUS_ADR_I[15] ), .SP(w_clk_cpu_enable_339), 
            .CK(w_clk_cpu), .Q(sram_adr_c_15)) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_addr_i16.GSR = "ENABLED";
    PFUMX sram_addr_nxt_18__I_0_i1 (.BLUT(sram_addr_nxt_18__N_3187), .ALUT(\SHAREDBUS_ADR_I[0] ), 
          .C0(sram_addr_nxt_18__N_3069), .Z(sram_addr_nxt[0])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;
    FD1P3AX sram_addr_i15 (.D(\SHAREDBUS_ADR_I[14] ), .SP(w_clk_cpu_enable_339), 
            .CK(w_clk_cpu), .Q(sram_adr_c_14)) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_addr_i15.GSR = "ENABLED";
    FD1P3AX sram_addr_i14 (.D(n41435), .SP(w_clk_cpu_enable_339), .CK(w_clk_cpu), 
            .Q(sram_adr_c_13)) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_addr_i14.GSR = "ENABLED";
    LUT4 sram_addr_nxt_18__I_0_i2_4_lut (.A(n41478), .B(\LM32D_ADR_O[1] ), 
         .C(n26018), .D(n41412), .Z(sram_addr_nxt[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(333[8] 344[36])
    defparam sram_addr_nxt_18__I_0_i2_4_lut.init = 16'hca0a;
    FD1P3AX sram_addr_i13 (.D(\SHAREDBUS_ADR_I[12] ), .SP(w_clk_cpu_enable_339), 
            .CK(w_clk_cpu), .Q(sram_adr_c_12)) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_addr_i13.GSR = "ENABLED";
    FD1P3AX sram_addr_i12 (.D(\SHAREDBUS_ADR_I[11] ), .SP(w_clk_cpu_enable_339), 
            .CK(w_clk_cpu), .Q(sram_adr_c_11)) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_addr_i12.GSR = "ENABLED";
    LUT4 i23378_2_lut (.A(n41405), .B(sram_addr_nxt_18__N_3069), .Z(n26018)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i23378_2_lut.init = 16'heeee;
    FD1P3AX sram_addr_i11 (.D(\SHAREDBUS_ADR_I[10] ), .SP(w_clk_cpu_enable_339), 
            .CK(w_clk_cpu), .Q(sram_adr_c_10)) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_addr_i11.GSR = "ENABLED";
    FD1P3AX sram_addr_i10 (.D(\SHAREDBUS_ADR_I[9] ), .SP(w_clk_cpu_enable_339), 
            .CK(w_clk_cpu), .Q(sram_adr_c_9)) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_addr_i10.GSR = "ENABLED";
    PFUMX cycle_counter_nxt_1__I_0_i2 (.BLUT(cycle_counter_nxt_1__N_3177[1]), 
          .ALUT(acycle[1]), .C0(n41353), .Z(cycle_counter_nxt[1])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;
    FD1P3AX sram_addr_i9 (.D(\SHAREDBUS_ADR_I[8] ), .SP(w_clk_cpu_enable_339), 
            .CK(w_clk_cpu), .Q(sram_adr_c_8)) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_addr_i9.GSR = "ENABLED";
    FD1P3AX sram_addr_i8 (.D(\SHAREDBUS_ADR_I[7] ), .SP(w_clk_cpu_enable_339), 
            .CK(w_clk_cpu), .Q(sram_adr_c_7)) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_addr_i8.GSR = "ENABLED";
    FD1P3AX sram_addr_i7 (.D(\SHAREDBUS_ADR_I[6] ), .SP(w_clk_cpu_enable_339), 
            .CK(w_clk_cpu), .Q(sram_adr_c_6)) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_addr_i7.GSR = "ENABLED";
    FD1P3AX sram_addr_i6 (.D(\SHAREDBUS_ADR_I[5] ), .SP(w_clk_cpu_enable_339), 
            .CK(w_clk_cpu), .Q(sram_adr_c_5)) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_addr_i6.GSR = "ENABLED";
    FD1P3AX sram_addr_i5 (.D(\SHAREDBUS_ADR_I[4] ), .SP(w_clk_cpu_enable_339), 
            .CK(w_clk_cpu), .Q(sram_adr_c_4)) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_addr_i5.GSR = "ENABLED";
    FD1P3AX sram_addr_i4 (.D(\SHAREDBUS_ADR_I[3] ), .SP(w_clk_cpu_enable_339), 
            .CK(w_clk_cpu), .Q(sram_adr_c_3)) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_addr_i4.GSR = "ENABLED";
    FD1P3AX sram_addr_i3 (.D(\SHAREDBUS_ADR_I[2] ), .SP(w_clk_cpu_enable_339), 
            .CK(w_clk_cpu), .Q(sram_adr_c_2)) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_addr_i3.GSR = "ENABLED";
    FD1P3AX sram_addr_i2 (.D(sram_addr_nxt[1]), .SP(w_clk_cpu_enable_339), 
            .CK(w_clk_cpu), .Q(sram_adr_c_1)) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_addr_i2.GSR = "ENABLED";
    FD1P3AX cycle_counter_i1 (.D(cycle_counter_nxt[1]), .SP(w_clk_cpu_enable_349), 
            .CK(w_clk_cpu), .Q(cycle[1])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(216[7:45])
    defparam cycle_counter_i1.GSR = "ENABLED";
    FD1P3IX dly_i3 (.D(n29457), .SP(tmp_dat_o_nxt_31__N_3127), .CD(n633), 
            .CK(w_clk_cpu), .Q(dly[3])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam dly_i3.GSR = "ENABLED";
    FD1P3IX dly_i2 (.D(n29460), .SP(tmp_dat_o_nxt_31__N_3127), .CD(n633), 
            .CK(w_clk_cpu), .Q(dly[2])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam dly_i2.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_337_4_lut_4_lut (.A(LM32D_SEL_O[2]), .B(selected[0]), 
         .C(selected[1]), .D(LM32D_SEL_O[3]), .Z(n41424)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C)+!B !(C (D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(549[17:33])
    defparam i1_2_lut_rep_337_4_lut_4_lut.init = 16'h3c2c;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut (.A(selected[0]), .B(selected[1]), 
         .C(n38761), .D(LM32D_SEL_O[3]), .Z(PIO_OUT_7__N_3327)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C (D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(535[12:28])
    defparam i1_2_lut_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h6020;
    FD1P3AX dly_i1 (.D(dly_nxt[1]), .SP(w_clk_cpu_enable_363), .CK(w_clk_cpu), 
            .Q(dly[1])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam dly_i1.GSR = "ENABLED";
    LUT4 tmp_dat_o_nxt_31__I_151_i1_4_lut (.A(sramsram_data_in[0]), .B(n467[0]), 
         .C(n41405), .D(n7), .Z(tmp_dat_o_nxt_31__N_3094[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i1_4_lut.init = 16'hca0a;
    LUT4 mux_199_i1_4_lut (.A(n21518[0]), .B(sramsram_data_in[0]), .C(n41393), 
         .D(n24342), .Z(n467[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(555[10] 562[17])
    defparam mux_199_i1_4_lut.init = 16'hca0a;
    LUT4 i2_4_lut (.A(n41423), .B(n41490), .C(LM32D_SEL_O[1]), .D(LM32D_SEL_O[0]), 
         .Z(n25515)) /* synthesis lut_function=(!((B+(C (D)+!C !(D)))+!A)) */ ;
    defparam i2_4_lut.init = 16'h0220;
    LUT4 i3_4_lut_adj_435 (.A(dly[1]), .B(dly[0]), .C(dly[2]), .D(dly[3]), 
         .Z(n25664)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam i3_4_lut_adj_435.init = 16'hfffb;
    LUT4 i3_4_lut_adj_436 (.A(n25664), .B(n42723), .C(w_clk_cpu_enable_303), 
         .D(n41488), .Z(dly_nxt_3__N_3169)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i3_4_lut_adj_436.init = 16'h0004;
    LUT4 cycle_counter_nxt_1__I_0_i1_4_lut (.A(cycle[0]), .B(n41363), .C(n41353), 
         .D(cycle_counter_nxt_1__N_3179), .Z(cycle_counter_nxt[0])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(206[10] 210[41])
    defparam cycle_counter_nxt_1__I_0_i1_4_lut.init = 16'hc5ca;
    LUT4 i22086_2_lut (.A(LM32D_SEL_O[2]), .B(LM32D_SEL_O[3]), .Z(n24709)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i22086_2_lut.init = 16'h6666;
    LUT4 i1_2_lut (.A(cycle_counter_nxt_1__N_3179), .B(sram_addr_nxt_18__N_3069), 
         .Z(w_clk_cpu_enable_339)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 sram_addr_nxt_18__I_121_4_lut (.A(n41501), .B(n41500), .C(n42723), 
         .D(n41356), .Z(sram_addr_nxt_18__N_3069)) /* synthesis lut_function=(!(A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(329[10] 330[77])
    defparam sram_addr_nxt_18__I_121_4_lut.init = 16'h5d55;
    LUT4 i1_4_lut_4_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_SEL_O[0]), 
         .D(LM32D_SEL_O[1]), .Z(n39016)) /* synthesis lut_function=(!(A (B)+!A !(B (C+(D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(559[5:12])
    defparam i1_4_lut_4_lut.init = 16'h6662;
    LUT4 i23406_3_lut (.A(LM32D_DAT_O[8]), .B(LM32D_DAT_O[0]), .C(sram_data_out_nxt_7__N_3086), 
         .Z(n26047)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(354[11] 362[42])
    defparam i23406_3_lut.init = 16'hcaca;
    LUT4 i20784_1_lut (.A(state[1]), .Z(w_clk_cpu_enable_184)) /* synthesis lut_function=(!(A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(333[13:31])
    defparam i20784_1_lut.init = 16'h5555;
    PFUMX i21209 (.BLUT(n36688), .ALUT(n183), .C0(state[1]), .Z(n23818));
    LUT4 i23404_3_lut (.A(LM32D_DAT_O[24]), .B(LM32D_DAT_O[16]), .C(n22230), 
         .Z(n26045)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(358[11] 362[42])
    defparam i23404_3_lut.init = 16'hcaca;
    LUT4 sram_data_out_nxt_7__I_124_4_lut (.A(n38998), .B(n41500), .C(n31536), 
         .D(n41497), .Z(sram_data_out_nxt_7__N_3086)) /* synthesis lut_function=(!(A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(347[10] 348[95])
    defparam sram_data_out_nxt_7__I_124_4_lut.init = 16'h5d55;
    LUT4 i38025_2_lut (.A(sram_data_out_nxt_7__N_3086), .B(sram_data_out_nxt_7__N_3201), 
         .Z(n39339)) /* synthesis lut_function=(A+(B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(350[11] 362[42])
    defparam i38025_2_lut.init = 16'heeee;
    LUT4 i2_4_lut_adj_437 (.A(n41500), .B(sram_data_out_nxt_7__N_3203), 
         .C(n41374), .D(n37005), .Z(sram_data_out_nxt_7__N_3201)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(350[15] 352[69])
    defparam i2_4_lut_adj_437.init = 16'hffec;
    LUT4 i3_4_lut_adj_438 (.A(n5_adj_3938), .B(sram_data_out_nxt_7__N_3086), 
         .C(n39018), .D(n40734), .Z(w_clk_cpu_enable_900)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam i3_4_lut_adj_438.init = 16'hffef;
    LUT4 i1_2_lut_adj_439 (.A(sram_data_out_nxt_7__N_3201), .B(n22230), 
         .Z(n5_adj_3938)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_439.init = 16'heeee;
    LUT4 i1_2_lut_rep_409 (.A(cycle[0]), .B(cycle[1]), .Z(n41496)) /* synthesis lut_function=(!(A+!(B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(216[7:45])
    defparam i1_2_lut_rep_409.init = 16'h4444;
    LUT4 i1_2_lut_3_lut (.A(cycle[0]), .B(cycle[1]), .C(sramsram_data_in[1]), 
         .Z(n14)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(216[7:45])
    defparam i1_2_lut_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_3_lut_adj_440 (.A(cycle[0]), .B(cycle[1]), .C(sramsram_data_in[0]), 
         .Z(tmp_dat_o_nxt_31__N_3239[16])) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(216[7:45])
    defparam i1_2_lut_3_lut_adj_440.init = 16'h4040;
    LUT4 i1_2_lut_rep_287_2_lut_3_lut (.A(cycle[0]), .B(cycle[1]), .C(n41405), 
         .Z(n41374)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(216[7:45])
    defparam i1_2_lut_rep_287_2_lut_3_lut.init = 16'h0404;
    LUT4 i29675_2_lut_3_lut_3_lut_4_lut_3_lut (.A(cycle[0]), .B(cycle[1]), 
         .C(n41405), .Z(sram_addr_nxt_18__N_3187)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(216[7:45])
    defparam i29675_2_lut_3_lut_3_lut_4_lut_3_lut.init = 16'hfbfb;
    LUT4 i1_2_lut_rep_410 (.A(cycle[0]), .B(cycle[1]), .Z(n41497)) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(216[7:45])
    defparam i1_2_lut_rep_410.init = 16'h2222;
    LUT4 i22562_2_lut_3_lut_2_lut (.A(cycle[0]), .B(cycle[1]), .Z(cycle_counter_nxt_1__N_3177[1])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(216[7:45])
    defparam i22562_2_lut_3_lut_2_lut.init = 16'h9999;
    FD1P3AX tmp_dat_o_i0_i31 (.D(tmp_dat_o_nxt_31__N_3094[31]), .SP(w_clk_cpu_enable_527), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[31])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i31.GSR = "ENABLED";
    PFUMX state_1__I_0_260_Mux_0_i1 (.BLUT(state_nxt_1__N_3154), .ALUT(n38992), 
          .C0(state[0]), .Z(n1)) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;
    FD1P3AX tmp_dat_o_i0_i30 (.D(tmp_dat_o_nxt_31__N_3094[30]), .SP(w_clk_cpu_enable_527), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[30])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i30.GSR = "ENABLED";
    FD1P3AX tmp_dat_o_i0_i29 (.D(tmp_dat_o_nxt_31__N_3094[29]), .SP(w_clk_cpu_enable_527), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[29])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i29.GSR = "ENABLED";
    FD1P3AX tmp_dat_o_i0_i28 (.D(tmp_dat_o_nxt_31__N_3094[28]), .SP(w_clk_cpu_enable_527), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[28])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i28.GSR = "ENABLED";
    FD1P3AX tmp_dat_o_i0_i27 (.D(tmp_dat_o_nxt_31__N_3094[27]), .SP(w_clk_cpu_enable_527), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[27])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i27.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_448 (.A(cycle[0]), .B(cycle[1]), .Z(n42723)) /* synthesis lut_function=(A+(B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam i1_2_lut_rep_448.init = 16'heeee;
    FD1P3AX tmp_dat_o_i0_i26 (.D(tmp_dat_o_nxt_31__N_3094[26]), .SP(w_clk_cpu_enable_527), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[26])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i26.GSR = "ENABLED";
    FD1P3AX tmp_dat_o_i0_i25 (.D(tmp_dat_o_nxt_31__N_3094[25]), .SP(w_clk_cpu_enable_527), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[25])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i25.GSR = "ENABLED";
    FD1P3AX tmp_dat_o_i0_i24 (.D(tmp_dat_o_nxt_31__N_3094[24]), .SP(w_clk_cpu_enable_527), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[24])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i24.GSR = "ENABLED";
    FD1P3AX tmp_dat_o_i0_i23 (.D(tmp_dat_o_nxt_31__N_3094[23]), .SP(w_clk_cpu_enable_566), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[23])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i23.GSR = "ENABLED";
    FD1P3AX tmp_dat_o_i0_i22 (.D(tmp_dat_o_nxt_31__N_3094[22]), .SP(w_clk_cpu_enable_566), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[22])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i22.GSR = "ENABLED";
    LUT4 i21296_4_lut_else_3_lut (.A(n42723), .B(n25664), .C(state[1]), 
         .D(state[0]), .Z(n41618)) /* synthesis lut_function=(A (B (C (D))+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(206[14] 207[77])
    defparam i21296_4_lut_else_3_lut.init = 16'ha200;
    FD1P3AX tmp_dat_o_i0_i21 (.D(tmp_dat_o_nxt_31__N_3094[21]), .SP(w_clk_cpu_enable_566), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[21])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i21.GSR = "ENABLED";
    LUT4 i23439_3_lut (.A(LM32D_DAT_O[12]), .B(LM32D_DAT_O[4]), .C(sram_data_out_nxt_7__N_3086), 
         .Z(n26081)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(354[11] 362[42])
    defparam i23439_3_lut.init = 16'hcaca;
    LUT4 i23426_3_lut (.A(LM32D_DAT_O[28]), .B(LM32D_DAT_O[20]), .C(n22230), 
         .Z(n26067)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(358[11] 362[42])
    defparam i23426_3_lut.init = 16'hcaca;
    FD1P3AX tmp_dat_o_i0_i20 (.D(tmp_dat_o_nxt_31__N_3094[20]), .SP(w_clk_cpu_enable_566), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[20])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i20.GSR = "ENABLED";
    FD1P3AX tmp_dat_o_i0_i19 (.D(tmp_dat_o_nxt_31__N_3094[19]), .SP(w_clk_cpu_enable_566), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[19])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i19.GSR = "ENABLED";
    FD1P3AX tmp_dat_o_i0_i18 (.D(tmp_dat_o_nxt_31__N_3094[18]), .SP(w_clk_cpu_enable_566), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[18])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i18.GSR = "ENABLED";
    FD1P3AX tmp_dat_o_i0_i17 (.D(tmp_dat_o_nxt_31__N_3094[17]), .SP(w_clk_cpu_enable_577), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[17])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i17.GSR = "ENABLED";
    LUT4 i23465_3_lut (.A(LM32D_DAT_O[14]), .B(LM32D_DAT_O[6]), .C(sram_data_out_nxt_7__N_3086), 
         .Z(n26107)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(354[11] 362[42])
    defparam i23465_3_lut.init = 16'hcaca;
    FD1P3AX tmp_dat_o_i0_i16 (.D(tmp_dat_o_nxt_31__N_3094[16]), .SP(w_clk_cpu_enable_577), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[16])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i16.GSR = "ENABLED";
    FD1P3AX tmp_dat_o_i0_i15 (.D(tmp_dat_o_nxt_31__N_3094[15]), .SP(w_clk_cpu_enable_619), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[15])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i15.GSR = "ENABLED";
    LUT4 i3_4_lut_3_lut (.A(n41429), .B(n41393), .C(n41390), .Z(n28684)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i3_4_lut_3_lut.init = 16'h8080;
    FD1P3AX tmp_dat_o_i0_i14 (.D(tmp_dat_o_nxt_31__N_3094[14]), .SP(w_clk_cpu_enable_619), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[14])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i14.GSR = "ENABLED";
    FD1P3AX tmp_dat_o_i0_i13 (.D(tmp_dat_o_nxt_31__N_3094[13]), .SP(w_clk_cpu_enable_619), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[13])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i13.GSR = "ENABLED";
    FD1P3AX tmp_dat_o_i0_i12 (.D(tmp_dat_o_nxt_31__N_3094[12]), .SP(w_clk_cpu_enable_619), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[12])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i12.GSR = "ENABLED";
    FD1P3AX tmp_dat_o_i0_i11 (.D(tmp_dat_o_nxt_31__N_3094[11]), .SP(w_clk_cpu_enable_619), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[11])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i11.GSR = "ENABLED";
    FD1P3AX tmp_dat_o_i0_i10 (.D(tmp_dat_o_nxt_31__N_3094[10]), .SP(w_clk_cpu_enable_619), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[10])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i10.GSR = "ENABLED";
    FD1P3AX tmp_dat_o_i0_i9 (.D(tmp_dat_o_nxt_31__N_3094[9]), .SP(w_clk_cpu_enable_619), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[9])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i9.GSR = "ENABLED";
    FD1P3IX sram_data_out_i0 (.D(n26049), .SP(w_clk_cpu_enable_900), .CD(n26128), 
            .CK(w_clk_cpu), .Q(sramsram_data_out[0])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_data_out_i0.GSR = "ENABLED";
    FD1P3AX tmp_dat_o_i0_i8 (.D(tmp_dat_o_nxt_31__N_3094[8]), .SP(w_clk_cpu_enable_619), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[8])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i8.GSR = "ENABLED";
    FD1P3AX tmp_dat_o_i0_i7 (.D(tmp_dat_o_nxt_31__N_3094[7]), .SP(w_clk_cpu_enable_648), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[7])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i7.GSR = "ENABLED";
    FD1P3AX tmp_dat_o_i0_i6 (.D(tmp_dat_o_nxt_31__N_3094[6]), .SP(w_clk_cpu_enable_648), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[6])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i6.GSR = "ENABLED";
    LUT4 sram_addr_nxt_18__N_3073_bdd_4_lut_38226 (.A(n7_adj_99), .B(n7), 
         .C(n41405), .D(n41501), .Z(n40733)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A (B (C)))) */ ;
    defparam sram_addr_nxt_18__N_3073_bdd_4_lut_38226.init = 16'h153f;
    FD1P3AX tmp_dat_o_i0_i5 (.D(tmp_dat_o_nxt_31__N_3094[5]), .SP(w_clk_cpu_enable_648), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[5])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i5.GSR = "ENABLED";
    LUT4 i29426_2_lut_rep_413 (.A(state[0]), .B(state[1]), .Z(n41500)) /* synthesis lut_function=(A (B)) */ ;
    defparam i29426_2_lut_rep_413.init = 16'h8888;
    FD1P3AX tmp_dat_o_i0_i4 (.D(tmp_dat_o_nxt_31__N_3094[4]), .SP(w_clk_cpu_enable_648), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[4])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i4.GSR = "ENABLED";
    FD1P3AX tmp_dat_o_i0_i3 (.D(tmp_dat_o_nxt_31__N_3094[3]), .SP(w_clk_cpu_enable_648), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[3])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i3.GSR = "ENABLED";
    LUT4 b_c_bdd_2_lut_3_lut_4_lut (.A(state[0]), .B(state[1]), .C(n41341), 
         .D(cycle[0]), .Z(n41342)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam b_c_bdd_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i2_2_lut_rep_358_3_lut (.A(state[0]), .B(state[1]), .C(cycle[0]), 
         .Z(n41445)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_rep_358_3_lut.init = 16'h8080;
    LUT4 state_1__I_0_250_i3_2_lut_rep_414 (.A(state[0]), .B(state[1]), 
         .Z(n41501)) /* synthesis lut_function=(A+(B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(329[10:28])
    defparam state_1__I_0_250_i3_2_lut_rep_414.init = 16'heeee;
    FD1P3AX tmp_dat_o_i0_i2 (.D(tmp_dat_o_nxt_31__N_3094[2]), .SP(w_clk_cpu_enable_648), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[2])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i2.GSR = "ENABLED";
    FD1P3AX tmp_dat_o_i0_i1 (.D(tmp_dat_o_nxt_31__N_3094[1]), .SP(w_clk_cpu_enable_648), 
            .CK(w_clk_cpu), .Q(sramASRAM_DAT_O[1])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(606[7:37])
    defparam tmp_dat_o_i0_i1.GSR = "ENABLED";
    LUT4 i399_2_lut_3_lut_4_lut_3_lut (.A(state[0]), .B(state[1]), .C(dly_nxt_3__N_3169), 
         .Z(n633)) /* synthesis lut_function=(A (B+(C))+!A ((C)+!B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(329[10:28])
    defparam i399_2_lut_3_lut_4_lut_3_lut.init = 16'hf9f9;
    LUT4 i38096_2_lut_2_lut_3_lut_4_lut_2_lut_2_lut (.A(state[0]), .B(state[1]), 
         .Z(w_clk_cpu_enable_363)) /* synthesis lut_function=(A+!(B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(329[10:28])
    defparam i38096_2_lut_2_lut_3_lut_4_lut_2_lut_2_lut.init = 16'hbbbb;
    LUT4 i28978_2_lut_rep_366_3_lut_2_lut (.A(state[0]), .B(state[1]), .Z(n41453)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(329[10:28])
    defparam i28978_2_lut_rep_366_3_lut_2_lut.init = 16'h6666;
    LUT4 i2_3_lut_4_lut_4_lut (.A(n41390), .B(n7), .C(n41393), .D(n41392), 
         .Z(acycle[1])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(188[17] 192[16])
    defparam i2_3_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i23449_3_lut (.A(LM32D_DAT_O[30]), .B(LM32D_DAT_O[22]), .C(n22230), 
         .Z(n26091)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(358[11] 362[42])
    defparam i23449_3_lut.init = 16'hcaca;
    LUT4 i21296_4_lut_then_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(state[0]), 
         .D(state[1]), .Z(n41619)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam i21296_4_lut_then_3_lut_4_lut.init = 16'he000;
    LUT4 mux_19179_i12_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(sramsram_data_in[3]), 
         .D(sramASRAM_DAT_O[27]), .Z(n21518[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam mux_19179_i12_3_lut_4_lut.init = 16'hf1e0;
    LUT4 equal_19657_i7_2_lut_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(state[1]), 
         .D(state[0]), .Z(n7_adj_99)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam equal_19657_i7_2_lut_3_lut_4_lut.init = 16'hefff;
    PFUMX tmp_dat_o_nxt_31__I_151_i17 (.BLUT(tmp_dat_o_nxt_31__N_3239[16]), 
          .ALUT(tmp_dat_o_nxt_31__N_3207[16]), .C0(n41405), .Z(tmp_dat_o_nxt_31__N_3094[16])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;
    LUT4 i23467_3_lut (.A(LM32D_DAT_O[13]), .B(LM32D_DAT_O[5]), .C(sram_data_out_nxt_7__N_3086), 
         .Z(n26109)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(354[11] 362[42])
    defparam i23467_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_adj_441 (.A(cycle[0]), .B(cycle[1]), .C(n25664), 
         .Z(n38992)) /* synthesis lut_function=(A+(B+(C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam i1_2_lut_3_lut_adj_441.init = 16'hfefe;
    LUT4 mux_19179_i15_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(sramsram_data_in[6]), 
         .D(sramASRAM_DAT_O[30]), .Z(n21518[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam mux_19179_i15_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19179_i16_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(sramsram_data_in[7]), 
         .D(sramASRAM_DAT_O[31]), .Z(n21518[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam mux_19179_i16_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19179_i11_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(sramsram_data_in[2]), 
         .D(sramASRAM_DAT_O[26]), .Z(n21518[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam mux_19179_i11_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19179_i13_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(sramsram_data_in[4]), 
         .D(sramASRAM_DAT_O[28]), .Z(n21518[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam mux_19179_i13_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i23451_3_lut (.A(LM32D_DAT_O[29]), .B(LM32D_DAT_O[21]), .C(n22230), 
         .Z(n26093)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(358[11] 362[42])
    defparam i23451_3_lut.init = 16'hcaca;
    LUT4 mux_19179_i1_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(sramASRAM_DAT_O[16]), 
         .D(sramsram_data_in[0]), .Z(n21518[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam mux_19179_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19179_i5_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(sramASRAM_DAT_O[20]), 
         .D(sramsram_data_in[4]), .Z(n21518[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam mux_19179_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19179_i9_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(sramsram_data_in[0]), 
         .D(sramASRAM_DAT_O[24]), .Z(n21518[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam mux_19179_i9_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19179_i14_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(sramsram_data_in[5]), 
         .D(sramASRAM_DAT_O[29]), .Z(n21518[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam mux_19179_i14_3_lut_4_lut.init = 16'hf1e0;
    PFUMX i26834 (.BLUT(n14), .ALUT(tmp_dat_o_nxt_31__N_3207[17]), .C0(n41405), 
          .Z(tmp_dat_o_nxt_31__N_3094[17]));
    LUT4 mux_19179_i10_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(sramsram_data_in[1]), 
         .D(sramASRAM_DAT_O[25]), .Z(n21518[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam mux_19179_i10_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i23441_3_lut (.A(LM32D_DAT_O[11]), .B(LM32D_DAT_O[3]), .C(sram_data_out_nxt_7__N_3086), 
         .Z(n26083)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(354[11] 362[42])
    defparam i23441_3_lut.init = 16'hcaca;
    LUT4 mux_19179_i8_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(sramASRAM_DAT_O[23]), 
         .D(sramsram_data_in[7]), .Z(n21518[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam mux_19179_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i23428_3_lut (.A(LM32D_DAT_O[27]), .B(LM32D_DAT_O[19]), .C(n22230), 
         .Z(n26069)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(358[11] 362[42])
    defparam i23428_3_lut.init = 16'hcaca;
    LUT4 mux_19179_i7_3_lut_4_lut (.A(cycle[0]), .B(cycle[1]), .C(sramASRAM_DAT_O[22]), 
         .D(sramsram_data_in[6]), .Z(n21518[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam mux_19179_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i23443_3_lut (.A(LM32D_DAT_O[10]), .B(LM32D_DAT_O[2]), .C(sram_data_out_nxt_7__N_3086), 
         .Z(n26085)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(354[11] 362[42])
    defparam i23443_3_lut.init = 16'hcaca;
    LUT4 i23430_3_lut (.A(LM32D_DAT_O[26]), .B(LM32D_DAT_O[18]), .C(n22230), 
         .Z(n26071)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(358[11] 362[42])
    defparam i23430_3_lut.init = 16'hcaca;
    LUT4 i28940_4_lut (.A(dly[2]), .B(dly[3]), .C(dly[0]), .D(dly[1]), 
         .Z(n29457)) /* synthesis lut_function=(A (B)+!A (B (C+(D))+!B !(C+(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(108[21:24])
    defparam i28940_4_lut.init = 16'hccc9;
    LUT4 i26841_3_lut (.A(dly[0]), .B(dly[2]), .C(dly[1]), .Z(n29460)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(108[21:24])
    defparam i26841_3_lut.init = 16'hc9c9;
    LUT4 i23445_3_lut (.A(LM32D_DAT_O[9]), .B(LM32D_DAT_O[1]), .C(sram_data_out_nxt_7__N_3086), 
         .Z(n26087)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(354[11] 362[42])
    defparam i23445_3_lut.init = 16'hcaca;
    LUT4 i23432_3_lut (.A(LM32D_DAT_O[25]), .B(LM32D_DAT_O[17]), .C(n22230), 
         .Z(n26073)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(358[11] 362[42])
    defparam i23432_3_lut.init = 16'hcaca;
    LUT4 i23463_3_lut (.A(LM32D_DAT_O[15]), .B(LM32D_DAT_O[7]), .C(sram_data_out_nxt_7__N_3086), 
         .Z(n26105)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(354[11] 362[42])
    defparam i23463_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_adj_442 (.A(n41453), .B(dly_nxt_3__N_3169), .C(dly[0]), 
         .D(dly[1]), .Z(dly_nxt[1])) /* synthesis lut_function=((B+(C (D)+!C !(D)))+!A) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(151[7] 156[18])
    defparam i2_4_lut_adj_442.init = 16'hfddf;
    LUT4 i23447_3_lut (.A(LM32D_DAT_O[31]), .B(LM32D_DAT_O[23]), .C(n22230), 
         .Z(n26089)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(358[11] 362[42])
    defparam i23447_3_lut.init = 16'hcaca;
    LUT4 i38078_2_lut_3_lut_3_lut_4_lut (.A(n41488), .B(n25664), .C(n41496), 
         .D(n41405), .Z(w_clk_cpu_enable_577)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam i38078_2_lut_3_lut_3_lut_4_lut.init = 16'h1110;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n41488), .B(n25664), .C(n41405), .D(n41496), 
         .Z(w_clk_cpu_enable_566)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h1110;
    LUT4 i1_3_lut_3_lut_4_lut (.A(n41488), .B(n25664), .C(n41405), .D(n41478), 
         .Z(w_clk_cpu_enable_527)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam i1_3_lut_3_lut_4_lut.init = 16'h1011;
    LUT4 i38053_3_lut_3_lut_4_lut (.A(n41488), .B(n25664), .C(n42723), 
         .D(n41405), .Z(w_clk_cpu_enable_648)) /* synthesis lut_function=(!(A+(B+!((D)+!C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam i38053_3_lut_3_lut_4_lut.init = 16'h1101;
    LUT4 i1_3_lut_4_lut (.A(n41488), .B(n25664), .C(n41405), .D(n41497), 
         .Z(w_clk_cpu_enable_619)) /* synthesis lut_function=(!(A+(B+!(C+(D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(167[11] 170[9])
    defparam i1_3_lut_4_lut.init = 16'h1110;
    LUT4 i2_3_lut_3_lut_4_lut_4_lut (.A(n41479), .B(n41469), .C(n39016), 
         .D(n41455), .Z(n7)) /* synthesis lut_function=(A ((C)+!B)+!A ((C+!(D))+!B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(535[12:28])
    defparam i2_3_lut_3_lut_4_lut_4_lut.init = 16'hf3f7;
    LUT4 mux_9_i5_3_lut_4_lut_4_lut (.A(n41479), .B(\data[28] ), .C(\SHAREDBUS_DAT_I[28] ), 
         .D(n41455), .Z(n96[4])) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(535[12:28])
    defparam mux_9_i5_3_lut_4_lut_4_lut.init = 16'hf0e4;
    LUT4 mux_9_i6_3_lut_4_lut_4_lut (.A(n41479), .B(\data[29] ), .C(\SHAREDBUS_DAT_I[29] ), 
         .D(n41455), .Z(n96[5])) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(535[12:28])
    defparam mux_9_i6_3_lut_4_lut_4_lut.init = 16'hf0e4;
    LUT4 mux_9_i7_3_lut_4_lut_4_lut (.A(n41479), .B(\data[30] ), .C(\SHAREDBUS_DAT_I[30] ), 
         .D(n41455), .Z(n96[6])) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(535[12:28])
    defparam mux_9_i7_3_lut_4_lut_4_lut.init = 16'hf0e4;
    LUT4 mux_9_i8_3_lut_4_lut_4_lut (.A(n41479), .B(\data[31] ), .C(\SHAREDBUS_DAT_I[31] ), 
         .D(n41455), .Z(n96[7])) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(535[12:28])
    defparam mux_9_i8_3_lut_4_lut_4_lut.init = 16'hf0e4;
    LUT4 mux_9_i4_3_lut_4_lut_4_lut (.A(n41479), .B(\data[27] ), .C(\SHAREDBUS_DAT_I[27] ), 
         .D(n41455), .Z(n96[3])) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(535[12:28])
    defparam mux_9_i4_3_lut_4_lut_4_lut.init = 16'hf0e4;
    LUT4 mux_9_i3_3_lut_4_lut_4_lut (.A(n41479), .B(\data[26] ), .C(\SHAREDBUS_DAT_I[26] ), 
         .D(n41455), .Z(n96[2])) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(535[12:28])
    defparam mux_9_i3_3_lut_4_lut_4_lut.init = 16'hf0e4;
    LUT4 mux_9_i2_3_lut_4_lut_4_lut (.A(n41479), .B(\data[25] ), .C(\SHAREDBUS_DAT_I[25] ), 
         .D(n41455), .Z(n96[1])) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(535[12:28])
    defparam mux_9_i2_3_lut_4_lut_4_lut.init = 16'hf0e4;
    LUT4 mux_9_i1_3_lut_4_lut_4_lut (.A(n41479), .B(\data[24] ), .C(\SHAREDBUS_DAT_I[24] ), 
         .D(n41455), .Z(n96[0])) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(535[12:28])
    defparam mux_9_i1_3_lut_4_lut_4_lut.init = 16'hf0e4;
    LUT4 tmp_dat_o_nxt_31__I_151_i21_3_lut (.A(sramsram_data_in[4]), .B(tmp_dat_o_nxt_31__N_3207[20]), 
         .C(n41405), .Z(tmp_dat_o_nxt_31__N_3094[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i21_3_lut.init = 16'hcaca;
    LUT4 mux_200_i21_4_lut (.A(n21518[4]), .B(n28684), .C(n7), .D(sramsram_data_in[4]), 
         .Z(tmp_dat_o_nxt_31__N_3207[20])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(549[13] 562[17])
    defparam mux_200_i21_4_lut.init = 16'hca0a;
    LUT4 tmp_dat_o_nxt_31__I_151_i20_3_lut (.A(sramsram_data_in[3]), .B(\tmp_dat_o_nxt_31__N_3207[19] ), 
         .C(n41405), .Z(tmp_dat_o_nxt_31__N_3094[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i20_3_lut.init = 16'hcaca;
    LUT4 tmp_dat_o_nxt_31__I_151_i19_3_lut (.A(sramsram_data_in[2]), .B(tmp_dat_o_nxt_31__N_3207[18]), 
         .C(n41405), .Z(tmp_dat_o_nxt_31__N_3094[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i19_3_lut.init = 16'hcaca;
    FD1P3IX sram_data_out_i7 (.D(n26111), .SP(w_clk_cpu_enable_900), .CD(n26128), 
            .CK(w_clk_cpu), .Q(sramsram_data_out[7])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_data_out_i7.GSR = "ENABLED";
    LUT4 mux_200_i19_4_lut (.A(n21518[2]), .B(n28684), .C(n7), .D(sramsram_data_in[2]), 
         .Z(tmp_dat_o_nxt_31__N_3207[18])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(549[13] 562[17])
    defparam mux_200_i19_4_lut.init = 16'hca0a;
    LUT4 state_1__I_0_259_i3_2_lut_rep_401 (.A(state[0]), .B(state[1]), 
         .Z(n41488)) /* synthesis lut_function=((B)+!A) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(534[10:28])
    defparam state_1__I_0_259_i3_2_lut_rep_401.init = 16'hdddd;
    LUT4 i37900_2_lut_rep_391 (.A(cycle[0]), .B(cycle[1]), .Z(n41478)) /* synthesis lut_function=(!(A (B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(216[7:45])
    defparam i37900_2_lut_rep_391.init = 16'h7777;
    LUT4 i37789_2_lut_3_lut (.A(state[0]), .B(state[1]), .C(dly[0]), .Z(dly_nxt_3__N_3165[0])) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (C)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(534[10:28])
    defparam i37789_2_lut_3_lut.init = 16'hd2d2;
    LUT4 tmp_dat_o_nxt_31__I_151_i16_4_lut (.A(sramsram_data_in[7]), .B(n467[15]), 
         .C(n41405), .D(n7), .Z(tmp_dat_o_nxt_31__N_3094[15])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i16_4_lut.init = 16'hca0a;
    LUT4 state_1__I_0_259_i4_1_lut_2_lut (.A(state[0]), .B(state[1]), .Z(tmp_dat_o_nxt_31__N_3127)) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(534[10:28])
    defparam state_1__I_0_259_i4_1_lut_2_lut.init = 16'h2222;
    LUT4 i28971_2_lut_3_lut_4_lut (.A(state[0]), .B(state[1]), .C(n41490), 
         .D(LM32D_WE_O), .Z(sram_oen_c)) /* synthesis lut_function=((B+!(C+!(D)))+!A) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(534[10:28])
    defparam i28971_2_lut_3_lut_4_lut.init = 16'hdfdd;
    LUT4 mux_199_i16_4_lut (.A(n21518[15]), .B(sramsram_data_in[7]), .C(n41393), 
         .D(n36822), .Z(n467[15])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(555[10] 562[17])
    defparam mux_199_i16_4_lut.init = 16'h0aca;
    LUT4 tmp_dat_o_nxt_31__I_151_i32_3_lut (.A(sramsram_data_in[7]), .B(tmp_dat_o_nxt_31__N_3207[31]), 
         .C(n41405), .Z(tmp_dat_o_nxt_31__N_3094[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i32_3_lut.init = 16'hcaca;
    LUT4 mux_200_i32_4_lut (.A(n21518[15]), .B(sramsram_data_in[7]), .C(n7), 
         .D(n36806), .Z(tmp_dat_o_nxt_31__N_3207[31])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(549[13] 562[17])
    defparam mux_200_i32_4_lut.init = 16'h0aca;
    LUT4 i3_4_lut_adj_443 (.A(n41429), .B(n41393), .C(n41390), .D(n25515), 
         .Z(n36806)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(555[10] 562[17])
    defparam i3_4_lut_adj_443.init = 16'hffbf;
    LUT4 tmp_dat_o_nxt_31__I_151_i31_3_lut (.A(sramsram_data_in[6]), .B(tmp_dat_o_nxt_31__N_3207[30]), 
         .C(n41405), .Z(tmp_dat_o_nxt_31__N_3094[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i31_3_lut.init = 16'hcaca;
    LUT4 mux_200_i31_4_lut (.A(n21518[14]), .B(sramsram_data_in[6]), .C(n7), 
         .D(n36806), .Z(tmp_dat_o_nxt_31__N_3207[30])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(549[13] 562[17])
    defparam mux_200_i31_4_lut.init = 16'h0aca;
    LUT4 WBS_SEL_I_3__N_244_3__bdd_4_lut (.A(n41455), .B(n41479), .C(LM32D_SEL_O[0]), 
         .D(cycle[1]), .Z(n41341)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (B (D))) */ ;
    defparam WBS_SEL_I_3__N_244_3__bdd_4_lut.init = 16'hec00;
    LUT4 tmp_dat_o_nxt_31__I_151_i30_3_lut (.A(sramsram_data_in[5]), .B(tmp_dat_o_nxt_31__N_3207[29]), 
         .C(n41405), .Z(tmp_dat_o_nxt_31__N_3094[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i30_3_lut.init = 16'hcaca;
    LUT4 mux_200_i30_4_lut (.A(n21518[13]), .B(sramsram_data_in[5]), .C(n7), 
         .D(n36806), .Z(tmp_dat_o_nxt_31__N_3207[29])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(549[13] 562[17])
    defparam mux_200_i30_4_lut.init = 16'h0aca;
    FD1P3IX sram_data_out_i6 (.D(n26113), .SP(w_clk_cpu_enable_900), .CD(n26128), 
            .CK(w_clk_cpu), .Q(sramsram_data_out[6])) /* synthesis LSE_LINE_FILE_ID=39, LSE_LCOL=4, LSE_RCOL=36, LSE_LLINE=109, LSE_RLINE=128 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(371[8] 375[6])
    defparam sram_data_out_i6.GSR = "ENABLED";
    LUT4 SHAREDBUS_SEL_I_3__bdd_4_lut (.A(n41423), .B(n41426), .C(n41445), 
         .D(cycle[1]), .Z(n41343)) /* synthesis lut_function=(A (B)+!A !(((D)+!C)+!B)) */ ;
    defparam SHAREDBUS_SEL_I_3__bdd_4_lut.init = 16'h88c8;
    LUT4 tmp_dat_o_nxt_31__I_151_i29_3_lut (.A(sramsram_data_in[4]), .B(tmp_dat_o_nxt_31__N_3207[28]), 
         .C(n41405), .Z(tmp_dat_o_nxt_31__N_3094[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i29_3_lut.init = 16'hcaca;
    LUT4 mux_200_i29_4_lut (.A(n21518[12]), .B(sramsram_data_in[4]), .C(n7), 
         .D(n36806), .Z(tmp_dat_o_nxt_31__N_3207[28])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(549[13] 562[17])
    defparam mux_200_i29_4_lut.init = 16'h0aca;
    LUT4 tmp_dat_o_nxt_31__I_151_i28_3_lut (.A(sramsram_data_in[3]), .B(tmp_dat_o_nxt_31__N_3207[27]), 
         .C(n41405), .Z(tmp_dat_o_nxt_31__N_3094[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i28_3_lut.init = 16'hcaca;
    LUT4 mux_200_i28_4_lut (.A(n21518[11]), .B(sramsram_data_in[3]), .C(n7), 
         .D(n36806), .Z(tmp_dat_o_nxt_31__N_3207[27])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(549[13] 562[17])
    defparam mux_200_i28_4_lut.init = 16'h0aca;
    LUT4 tmp_dat_o_nxt_31__I_151_i27_3_lut (.A(sramsram_data_in[2]), .B(tmp_dat_o_nxt_31__N_3207[26]), 
         .C(n41405), .Z(tmp_dat_o_nxt_31__N_3094[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i27_3_lut.init = 16'hcaca;
    LUT4 mux_200_i27_4_lut (.A(n21518[10]), .B(sramsram_data_in[2]), .C(n7), 
         .D(n36806), .Z(tmp_dat_o_nxt_31__N_3207[26])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(549[13] 562[17])
    defparam mux_200_i27_4_lut.init = 16'h0aca;
    LUT4 tmp_dat_o_nxt_31__I_151_i26_3_lut (.A(sramsram_data_in[1]), .B(tmp_dat_o_nxt_31__N_3207[25]), 
         .C(n41405), .Z(tmp_dat_o_nxt_31__N_3094[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i26_3_lut.init = 16'hcaca;
    LUT4 mux_200_i26_4_lut (.A(n21518[9]), .B(sramsram_data_in[1]), .C(n7), 
         .D(n36806), .Z(tmp_dat_o_nxt_31__N_3207[25])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(549[13] 562[17])
    defparam mux_200_i26_4_lut.init = 16'h0aca;
    LUT4 tmp_dat_o_nxt_31__I_151_i25_3_lut (.A(sramsram_data_in[0]), .B(tmp_dat_o_nxt_31__N_3207[24]), 
         .C(n41405), .Z(tmp_dat_o_nxt_31__N_3094[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i25_3_lut.init = 16'hcaca;
    LUT4 mux_200_i25_4_lut (.A(n21518[8]), .B(sramsram_data_in[0]), .C(n7), 
         .D(n36806), .Z(tmp_dat_o_nxt_31__N_3207[24])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(549[13] 562[17])
    defparam mux_200_i25_4_lut.init = 16'h0aca;
    LUT4 tmp_dat_o_nxt_31__I_151_i24_3_lut (.A(sramsram_data_in[7]), .B(tmp_dat_o_nxt_31__N_3207[23]), 
         .C(n41405), .Z(tmp_dat_o_nxt_31__N_3094[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i24_3_lut.init = 16'hcaca;
    LUT4 mux_200_i24_4_lut (.A(n21518[7]), .B(n28684), .C(n7), .D(sramsram_data_in[7]), 
         .Z(tmp_dat_o_nxt_31__N_3207[23])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(549[13] 562[17])
    defparam mux_200_i24_4_lut.init = 16'hca0a;
    LUT4 tmp_dat_o_nxt_31__I_151_i23_3_lut (.A(sramsram_data_in[6]), .B(tmp_dat_o_nxt_31__N_3207[22]), 
         .C(n41405), .Z(tmp_dat_o_nxt_31__N_3094[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i23_3_lut.init = 16'hcaca;
    LUT4 mux_200_i23_4_lut (.A(n21518[6]), .B(n28684), .C(n7), .D(sramsram_data_in[6]), 
         .Z(tmp_dat_o_nxt_31__N_3207[22])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(549[13] 562[17])
    defparam mux_200_i23_4_lut.init = 16'hca0a;
    PFUMX i38623 (.BLUT(n41618), .ALUT(n41619), .C0(w_clk_cpu_enable_303), 
          .Z(cycle_counter_nxt_1__N_3179));
    LUT4 tmp_dat_o_nxt_31__I_151_i22_3_lut (.A(sramsram_data_in[5]), .B(tmp_dat_o_nxt_31__N_3207[21]), 
         .C(n41405), .Z(tmp_dat_o_nxt_31__N_3094[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(544[13] 562[17])
    defparam tmp_dat_o_nxt_31__I_151_i22_3_lut.init = 16'hcaca;
    LUT4 mux_200_i22_4_lut (.A(n21518[5]), .B(n28684), .C(n7), .D(sramsram_data_in[5]), 
         .Z(tmp_dat_o_nxt_31__N_3207[21])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/asram_top/rtl/verilog/asram_core.v(549[13] 562[17])
    defparam mux_200_i22_4_lut.init = 16'hca0a;
    
endmodule
//
// Verilog Description of module \gpio(DATA_WIDTH=32'b0100000,INPUT_WIDTH=32'b01,OUTPUT_WIDTH=32'b01,EDGE=1,POSE_EDGE_IRQ=1,INPUT_PORTS_ONLY=0,OUTPUT_PORTS_ONLY=1) 
//

module \gpio(DATA_WIDTH=32'b0100000,INPUT_WIDTH=32'b01,OUTPUT_WIDTH=32'b01,EDGE=1,POSE_EDGE_IRQ=1,INPUT_PORTS_ONLY=0,OUTPUT_PORTS_ONLY=1)  (gpioGPIO_ACK_O, 
            n93, n41366, w_clk_cpu, \counter[0] , PIO_OUT_7__N_3327, 
            \SHAREDBUS_DAT_I[24] , \counter[1] , \SHAREDBUS_DAT_I[25] , 
            \counter[2] , \SHAREDBUS_DAT_I[26] , w_clk_cpu_enable_303, 
            \SHAREDBUS_ADR_I[2] , \SHAREDBUS_ADR_I[3] , n38761, \counter[4] , 
            \SHAREDBUS_DAT_I[28] , \counter[5] , \SHAREDBUS_DAT_I[29] , 
            \counter[6] , \SHAREDBUS_DAT_I[30] , \counter[7] , \SHAREDBUS_DAT_I[31] , 
            \counter[8] , PIO_OUT_15__N_3318, \SHAREDBUS_DAT_I[16] , \counter[9] , 
            \SHAREDBUS_DAT_I[17] , \counter[10] , \SHAREDBUS_DAT_I[18] , 
            \counter[11] , \SHAREDBUS_DAT_I[19] , \counter[12] , \SHAREDBUS_DAT_I[20] , 
            \counter[13] , \SHAREDBUS_DAT_I[21] , \counter[14] , \SHAREDBUS_DAT_I[22] , 
            \counter[15] , \SHAREDBUS_DAT_I[23] , \counter[3] , \SHAREDBUS_DAT_I[27] ) /* synthesis syn_module_defined=1 */ ;
    output gpioGPIO_ACK_O;
    input [0:0]n93;
    input n41366;
    input w_clk_cpu;
    output \counter[0] ;
    input PIO_OUT_7__N_3327;
    input \SHAREDBUS_DAT_I[24] ;
    output \counter[1] ;
    input \SHAREDBUS_DAT_I[25] ;
    output \counter[2] ;
    input \SHAREDBUS_DAT_I[26] ;
    input w_clk_cpu_enable_303;
    input \SHAREDBUS_ADR_I[2] ;
    input \SHAREDBUS_ADR_I[3] ;
    output n38761;
    output \counter[4] ;
    input \SHAREDBUS_DAT_I[28] ;
    output \counter[5] ;
    input \SHAREDBUS_DAT_I[29] ;
    output \counter[6] ;
    input \SHAREDBUS_DAT_I[30] ;
    output \counter[7] ;
    input \SHAREDBUS_DAT_I[31] ;
    output \counter[8] ;
    input PIO_OUT_15__N_3318;
    input \SHAREDBUS_DAT_I[16] ;
    output \counter[9] ;
    input \SHAREDBUS_DAT_I[17] ;
    output \counter[10] ;
    input \SHAREDBUS_DAT_I[18] ;
    output \counter[11] ;
    input \SHAREDBUS_DAT_I[19] ;
    output \counter[12] ;
    input \SHAREDBUS_DAT_I[20] ;
    output \counter[13] ;
    input \SHAREDBUS_DAT_I[21] ;
    output \counter[14] ;
    input \SHAREDBUS_DAT_I[22] ;
    output \counter[15] ;
    input \SHAREDBUS_DAT_I[23] ;
    output \counter[3] ;
    input \SHAREDBUS_DAT_I[27] ;
    
    wire w_clk_cpu /* synthesis SET_AS_NETWORK=w_clk_cpu, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(22[6:15])
    
    wire PIO_OUT_31__N_3298;
    
    LUT4 i2_3_lut (.A(gpioGPIO_ACK_O), .B(n93[0]), .C(n41366), .Z(PIO_OUT_31__N_3298)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/gpio/rtl/verilog/gpio.v(188[14:48])
    defparam i2_3_lut.init = 16'h4040;
    FD1S3AX GPIO_ACK_O_469 (.D(PIO_OUT_31__N_3298), .CK(w_clk_cpu), .Q(gpioGPIO_ACK_O)) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=34, LSE_LLINE=623, LSE_RLINE=639 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/gpio/rtl/verilog/gpio.v(188[11] 191[33])
    defparam GPIO_ACK_O_469.GSR = "ENABLED";
    FD1P3AX PIO_DATA_0__470 (.D(\SHAREDBUS_DAT_I[24] ), .SP(PIO_OUT_7__N_3327), 
            .CK(w_clk_cpu), .Q(\counter[0] ));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/gpio/rtl/verilog/gpio.v(258[11] 259[62])
    defparam PIO_DATA_0__470.GSR = "ENABLED";
    FD1P3AX PIO_DATA_1__471 (.D(\SHAREDBUS_DAT_I[25] ), .SP(PIO_OUT_7__N_3327), 
            .CK(w_clk_cpu), .Q(\counter[1] ));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/gpio/rtl/verilog/gpio.v(258[11] 259[62])
    defparam PIO_DATA_1__471.GSR = "ENABLED";
    FD1P3AX PIO_DATA_2__472 (.D(\SHAREDBUS_DAT_I[26] ), .SP(PIO_OUT_7__N_3327), 
            .CK(w_clk_cpu), .Q(\counter[2] ));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/gpio/rtl/verilog/gpio.v(258[11] 259[62])
    defparam PIO_DATA_2__472.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(PIO_OUT_31__N_3298), .B(w_clk_cpu_enable_303), .C(\SHAREDBUS_ADR_I[2] ), 
         .D(\SHAREDBUS_ADR_I[3] ), .Z(n38761)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/gpio/rtl/verilog/gpio.v(188[14:48])
    defparam i2_4_lut.init = 16'h0008;
    FD1P3AX PIO_DATA_4__474 (.D(\SHAREDBUS_DAT_I[28] ), .SP(PIO_OUT_7__N_3327), 
            .CK(w_clk_cpu), .Q(\counter[4] ));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/gpio/rtl/verilog/gpio.v(258[11] 259[62])
    defparam PIO_DATA_4__474.GSR = "ENABLED";
    FD1P3AX PIO_DATA_5__475 (.D(\SHAREDBUS_DAT_I[29] ), .SP(PIO_OUT_7__N_3327), 
            .CK(w_clk_cpu), .Q(\counter[5] ));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/gpio/rtl/verilog/gpio.v(258[11] 259[62])
    defparam PIO_DATA_5__475.GSR = "ENABLED";
    FD1P3AX PIO_DATA_6__476 (.D(\SHAREDBUS_DAT_I[30] ), .SP(PIO_OUT_7__N_3327), 
            .CK(w_clk_cpu), .Q(\counter[6] ));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/gpio/rtl/verilog/gpio.v(258[11] 259[62])
    defparam PIO_DATA_6__476.GSR = "ENABLED";
    FD1P3AX PIO_DATA_7__477 (.D(\SHAREDBUS_DAT_I[31] ), .SP(PIO_OUT_7__N_3327), 
            .CK(w_clk_cpu), .Q(\counter[7] ));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/gpio/rtl/verilog/gpio.v(258[11] 259[62])
    defparam PIO_DATA_7__477.GSR = "ENABLED";
    FD1P3AX PIO_DATA_8__478 (.D(\SHAREDBUS_DAT_I[16] ), .SP(PIO_OUT_15__N_3318), 
            .CK(w_clk_cpu), .Q(\counter[8] ));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/gpio/rtl/verilog/gpio.v(268[14] 269[58])
    defparam PIO_DATA_8__478.GSR = "ENABLED";
    FD1P3AX PIO_DATA_9__479 (.D(\SHAREDBUS_DAT_I[17] ), .SP(PIO_OUT_15__N_3318), 
            .CK(w_clk_cpu), .Q(\counter[9] ));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/gpio/rtl/verilog/gpio.v(268[14] 269[58])
    defparam PIO_DATA_9__479.GSR = "ENABLED";
    FD1P3AX PIO_DATA_10__480 (.D(\SHAREDBUS_DAT_I[18] ), .SP(PIO_OUT_15__N_3318), 
            .CK(w_clk_cpu), .Q(\counter[10] ));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/gpio/rtl/verilog/gpio.v(268[14] 269[58])
    defparam PIO_DATA_10__480.GSR = "ENABLED";
    FD1P3AX PIO_DATA_11__481 (.D(\SHAREDBUS_DAT_I[19] ), .SP(PIO_OUT_15__N_3318), 
            .CK(w_clk_cpu), .Q(\counter[11] ));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/gpio/rtl/verilog/gpio.v(268[14] 269[58])
    defparam PIO_DATA_11__481.GSR = "ENABLED";
    FD1P3AX PIO_DATA_12__482 (.D(\SHAREDBUS_DAT_I[20] ), .SP(PIO_OUT_15__N_3318), 
            .CK(w_clk_cpu), .Q(\counter[12] ));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/gpio/rtl/verilog/gpio.v(268[14] 269[58])
    defparam PIO_DATA_12__482.GSR = "ENABLED";
    FD1P3AX PIO_DATA_13__483 (.D(\SHAREDBUS_DAT_I[21] ), .SP(PIO_OUT_15__N_3318), 
            .CK(w_clk_cpu), .Q(\counter[13] ));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/gpio/rtl/verilog/gpio.v(268[14] 269[58])
    defparam PIO_DATA_13__483.GSR = "ENABLED";
    FD1P3AX PIO_DATA_14__484 (.D(\SHAREDBUS_DAT_I[22] ), .SP(PIO_OUT_15__N_3318), 
            .CK(w_clk_cpu), .Q(\counter[14] ));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/gpio/rtl/verilog/gpio.v(268[14] 269[58])
    defparam PIO_DATA_14__484.GSR = "ENABLED";
    FD1P3AX PIO_DATA_15__485 (.D(\SHAREDBUS_DAT_I[23] ), .SP(PIO_OUT_15__N_3318), 
            .CK(w_clk_cpu), .Q(\counter[15] ));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/gpio/rtl/verilog/gpio.v(268[14] 269[58])
    defparam PIO_DATA_15__485.GSR = "ENABLED";
    FD1P3AX PIO_DATA_3__473 (.D(\SHAREDBUS_DAT_I[27] ), .SP(PIO_OUT_7__N_3327), 
            .CK(w_clk_cpu), .Q(\counter[3] ));   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/gpio/rtl/verilog/gpio.v(258[11] 259[62])
    defparam PIO_DATA_3__473.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module arbiter2
//

module arbiter2 (n41426, n41405, n41424, n31536, selected, \selected_1__N_344[0] , 
            w_clk_cpu, LM32D_SEL_O, LM32D_WE_O, w_clk_cpu_enable_303, 
            n92, n39983, \LM32I_ADR_O[11] , \LM32D_ADR_O[11] , \SHAREDBUS_ADR_I[11] , 
            n25515, n41392, n38761, PIO_OUT_15__N_3318, n41344, n22230, 
            \LM32I_ADR_O[5] , \LM32D_ADR_O[5] , \SHAREDBUS_ADR_I[5] , 
            \LM32I_ADR_O[8] , \LM32D_ADR_O[8] , \SHAREDBUS_ADR_I[8] , 
            \LM32I_ADR_O[12] , \LM32D_ADR_O[12] , \SHAREDBUS_ADR_I[12] , 
            w_clk_cpu_enable_900, n26128, \LM32I_ADR_O[17] , \LM32D_ADR_O[17] , 
            \SHAREDBUS_ADR_I[17] , \LM32I_ADR_O[16] , \LM32D_ADR_O[16] , 
            \SHAREDBUS_ADR_I[16] , \LM32I_ADR_O[18] , \LM32D_ADR_O[18] , 
            \SHAREDBUS_ADR_I[18] , \LM32I_ADR_O[15] , \LM32D_ADR_O[15] , 
            \SHAREDBUS_ADR_I[15] , \LM32I_ADR_O[14] , \LM32D_ADR_O[14] , 
            \SHAREDBUS_ADR_I[14] , \LM32D_DAT_O[24] , \SHAREDBUS_DAT_I[24] , 
            \LM32D_DAT_O[25] , \SHAREDBUS_DAT_I[25] , \SHAREDBUS_SEL_I[1] , 
            n41429, \LM32I_ADR_O[19] , \LM32D_ADR_O[19] , \SHAREDBUS_ADR_I[19] , 
            \LM32I_ADR_O[7] , \LM32D_ADR_O[7] , \SHAREDBUS_ADR_I[7] , 
            \LM32I_ADR_O[10] , \LM32D_ADR_O[10] , \SHAREDBUS_ADR_I[10] , 
            \LM32I_ADR_O[9] , \LM32D_ADR_O[9] , \SHAREDBUS_ADR_I[9] , 
            \LM32I_ADR_O[6] , \LM32D_ADR_O[6] , \SHAREDBUS_ADR_I[6] , 
            \LM32I_ADR_O[4] , \LM32D_ADR_O[4] , \SHAREDBUS_ADR_I[4] , 
            \LM32I_ADR_O[31] , \LM32D_ADR_O[31] , n41442, n41423, \LM32I_ADR_O[13] , 
            \LM32D_ADR_O[13] , n41435, \LM32I_ADR_O[22] , \LM32D_ADR_O[22] , 
            \SHAREDBUS_ADR_I[22] , \LM32I_ADR_O[26] , \LM32D_ADR_O[26] , 
            \SHAREDBUS_ADR_I[26] , \LM32I_ADR_O[25] , \LM32D_ADR_O[25] , 
            \SHAREDBUS_ADR_I[25] , \LM32I_ADR_O[24] , \LM32D_ADR_O[24] , 
            \SHAREDBUS_ADR_I[24] , \LM32I_ADR_O[27] , \LM32D_ADR_O[27] , 
            \SHAREDBUS_ADR_I[27] , \LM32I_ADR_O[28] , \LM32D_ADR_O[28] , 
            \SHAREDBUS_ADR_I[28] , \LM32D_DAT_O[26] , \SHAREDBUS_DAT_I[26] , 
            \LM32D_DAT_O[28] , \SHAREDBUS_DAT_I[28] , \LM32I_ADR_O[29] , 
            \LM32D_ADR_O[29] , \SHAREDBUS_ADR_I[29] , \LM32D_DAT_O[29] , 
            \SHAREDBUS_DAT_I[29] , \LM32D_DAT_O[30] , \SHAREDBUS_DAT_I[30] , 
            \LM32D_DAT_O[31] , \SHAREDBUS_DAT_I[31] , \LM32D_DAT_O[18] , 
            \SHAREDBUS_DAT_I[18] , \LM32D_DAT_O[19] , \SHAREDBUS_DAT_I[19] , 
            \LM32I_ADR_O[23] , \LM32D_ADR_O[23] , \SHAREDBUS_ADR_I[23] , 
            \LM32I_ADR_O[30] , \LM32D_ADR_O[30] , \SHAREDBUS_ADR_I[30] , 
            \LM32D_DAT_O[20] , \SHAREDBUS_DAT_I[20] , \LM32I_ADR_O[21] , 
            \LM32D_ADR_O[21] , \SHAREDBUS_ADR_I[21] , \LM32I_ADR_O[2] , 
            \LM32D_ADR_O[2] , \SHAREDBUS_ADR_I[2] , \LM32D_DAT_O[21] , 
            \SHAREDBUS_DAT_I[21] , \LM32I_ADR_O[3] , \LM32D_ADR_O[3] , 
            \SHAREDBUS_ADR_I[3] , \LM32D_DAT_O[22] , \SHAREDBUS_DAT_I[22] , 
            \LM32D_DAT_O[23] , \SHAREDBUS_DAT_I[23] , \LM32D_DAT_O[27] , 
            \SHAREDBUS_DAT_I[27] , \LM32I_ADR_O[20] , \LM32D_ADR_O[20] , 
            \SHAREDBUS_ADR_I[20] , LM32I_CYC_O, LM32D_CYC_O, LM32D_STB_O, 
            n93, n41479, n38998, n41393, n41469, \data[19] , n87, 
            n41390, n41363, \SHAREDBUS_DAT_I[16] , \data[16] , \SHAREDBUS_DAT_I[17] , 
            \data[17] , \data[23] , \data[18] , \data[22] , \data[20] , 
            \data[21] , n41490, n24709, n41412, n41455, \LM32D_DAT_O[17] , 
            tmp_ack_o, \genblk5.tmp_ack_o_d , n41421, n42723, n25664, 
            n36688, n24342, n36822, n37005, \LM32D_DAT_O[16] , n41352, 
            n76, n39016, n39018, n21531, \sramsram_data_in[3] , n7, 
            n28684, \tmp_dat_o_nxt_31__N_3207[19] , n38871, bus_error_f_N_1764, 
            \LM32D_ADR_O[0] , \SHAREDBUS_ADR_I[0] ) /* synthesis syn_module_defined=1 */ ;
    output n41426;
    output n41405;
    input n41424;
    output n31536;
    output [1:0]selected;
    input \selected_1__N_344[0] ;
    input w_clk_cpu;
    input [3:0]LM32D_SEL_O;
    input LM32D_WE_O;
    output w_clk_cpu_enable_303;
    output [0:0]n92;
    output n39983;
    input \LM32I_ADR_O[11] ;
    input \LM32D_ADR_O[11] ;
    output \SHAREDBUS_ADR_I[11] ;
    input n25515;
    output n41392;
    input n38761;
    output PIO_OUT_15__N_3318;
    input n41344;
    output n22230;
    input \LM32I_ADR_O[5] ;
    input \LM32D_ADR_O[5] ;
    output \SHAREDBUS_ADR_I[5] ;
    input \LM32I_ADR_O[8] ;
    input \LM32D_ADR_O[8] ;
    output \SHAREDBUS_ADR_I[8] ;
    input \LM32I_ADR_O[12] ;
    input \LM32D_ADR_O[12] ;
    output \SHAREDBUS_ADR_I[12] ;
    input w_clk_cpu_enable_900;
    output n26128;
    input \LM32I_ADR_O[17] ;
    input \LM32D_ADR_O[17] ;
    output \SHAREDBUS_ADR_I[17] ;
    input \LM32I_ADR_O[16] ;
    input \LM32D_ADR_O[16] ;
    output \SHAREDBUS_ADR_I[16] ;
    input \LM32I_ADR_O[18] ;
    input \LM32D_ADR_O[18] ;
    output \SHAREDBUS_ADR_I[18] ;
    input \LM32I_ADR_O[15] ;
    input \LM32D_ADR_O[15] ;
    output \SHAREDBUS_ADR_I[15] ;
    input \LM32I_ADR_O[14] ;
    input \LM32D_ADR_O[14] ;
    output \SHAREDBUS_ADR_I[14] ;
    input \LM32D_DAT_O[24] ;
    output \SHAREDBUS_DAT_I[24] ;
    input \LM32D_DAT_O[25] ;
    output \SHAREDBUS_DAT_I[25] ;
    output \SHAREDBUS_SEL_I[1] ;
    output n41429;
    input \LM32I_ADR_O[19] ;
    input \LM32D_ADR_O[19] ;
    output \SHAREDBUS_ADR_I[19] ;
    input \LM32I_ADR_O[7] ;
    input \LM32D_ADR_O[7] ;
    output \SHAREDBUS_ADR_I[7] ;
    input \LM32I_ADR_O[10] ;
    input \LM32D_ADR_O[10] ;
    output \SHAREDBUS_ADR_I[10] ;
    input \LM32I_ADR_O[9] ;
    input \LM32D_ADR_O[9] ;
    output \SHAREDBUS_ADR_I[9] ;
    input \LM32I_ADR_O[6] ;
    input \LM32D_ADR_O[6] ;
    output \SHAREDBUS_ADR_I[6] ;
    input \LM32I_ADR_O[4] ;
    input \LM32D_ADR_O[4] ;
    output \SHAREDBUS_ADR_I[4] ;
    input \LM32I_ADR_O[31] ;
    input \LM32D_ADR_O[31] ;
    output n41442;
    output n41423;
    input \LM32I_ADR_O[13] ;
    input \LM32D_ADR_O[13] ;
    output n41435;
    input \LM32I_ADR_O[22] ;
    input \LM32D_ADR_O[22] ;
    output \SHAREDBUS_ADR_I[22] ;
    input \LM32I_ADR_O[26] ;
    input \LM32D_ADR_O[26] ;
    output \SHAREDBUS_ADR_I[26] ;
    input \LM32I_ADR_O[25] ;
    input \LM32D_ADR_O[25] ;
    output \SHAREDBUS_ADR_I[25] ;
    input \LM32I_ADR_O[24] ;
    input \LM32D_ADR_O[24] ;
    output \SHAREDBUS_ADR_I[24] ;
    input \LM32I_ADR_O[27] ;
    input \LM32D_ADR_O[27] ;
    output \SHAREDBUS_ADR_I[27] ;
    input \LM32I_ADR_O[28] ;
    input \LM32D_ADR_O[28] ;
    output \SHAREDBUS_ADR_I[28] ;
    input \LM32D_DAT_O[26] ;
    output \SHAREDBUS_DAT_I[26] ;
    input \LM32D_DAT_O[28] ;
    output \SHAREDBUS_DAT_I[28] ;
    input \LM32I_ADR_O[29] ;
    input \LM32D_ADR_O[29] ;
    output \SHAREDBUS_ADR_I[29] ;
    input \LM32D_DAT_O[29] ;
    output \SHAREDBUS_DAT_I[29] ;
    input \LM32D_DAT_O[30] ;
    output \SHAREDBUS_DAT_I[30] ;
    input \LM32D_DAT_O[31] ;
    output \SHAREDBUS_DAT_I[31] ;
    input \LM32D_DAT_O[18] ;
    output \SHAREDBUS_DAT_I[18] ;
    input \LM32D_DAT_O[19] ;
    output \SHAREDBUS_DAT_I[19] ;
    input \LM32I_ADR_O[23] ;
    input \LM32D_ADR_O[23] ;
    output \SHAREDBUS_ADR_I[23] ;
    input \LM32I_ADR_O[30] ;
    input \LM32D_ADR_O[30] ;
    output \SHAREDBUS_ADR_I[30] ;
    input \LM32D_DAT_O[20] ;
    output \SHAREDBUS_DAT_I[20] ;
    input \LM32I_ADR_O[21] ;
    input \LM32D_ADR_O[21] ;
    output \SHAREDBUS_ADR_I[21] ;
    input \LM32I_ADR_O[2] ;
    input \LM32D_ADR_O[2] ;
    output \SHAREDBUS_ADR_I[2] ;
    input \LM32D_DAT_O[21] ;
    output \SHAREDBUS_DAT_I[21] ;
    input \LM32I_ADR_O[3] ;
    input \LM32D_ADR_O[3] ;
    output \SHAREDBUS_ADR_I[3] ;
    input \LM32D_DAT_O[22] ;
    output \SHAREDBUS_DAT_I[22] ;
    input \LM32D_DAT_O[23] ;
    output \SHAREDBUS_DAT_I[23] ;
    input \LM32D_DAT_O[27] ;
    output \SHAREDBUS_DAT_I[27] ;
    input \LM32I_ADR_O[20] ;
    input \LM32D_ADR_O[20] ;
    output \SHAREDBUS_ADR_I[20] ;
    input LM32I_CYC_O;
    input LM32D_CYC_O;
    input LM32D_STB_O;
    output [0:0]n93;
    output n41479;
    output n38998;
    output n41393;
    output n41469;
    input \data[19] ;
    output [7:0]n87;
    output n41390;
    output n41363;
    output \SHAREDBUS_DAT_I[16] ;
    input \data[16] ;
    output \SHAREDBUS_DAT_I[17] ;
    input \data[17] ;
    input \data[23] ;
    input \data[18] ;
    input \data[22] ;
    input \data[20] ;
    input \data[21] ;
    output n41490;
    input n24709;
    output n41412;
    output n41455;
    input \LM32D_DAT_O[17] ;
    input tmp_ack_o;
    input \genblk5.tmp_ack_o_d ;
    output n41421;
    input n42723;
    input n25664;
    output n36688;
    output n24342;
    output n36822;
    output n37005;
    input \LM32D_DAT_O[16] ;
    input n41352;
    input [0:0]n76;
    input n39016;
    output n39018;
    input n21531;
    input \sramsram_data_in[3] ;
    input n7;
    input n28684;
    output \tmp_dat_o_nxt_31__N_3207[19] ;
    input n38871;
    output bus_error_f_N_1764;
    input \LM32D_ADR_O[0] ;
    output \SHAREDBUS_ADR_I[0] ;
    
    wire w_clk_cpu /* synthesis SET_AS_NETWORK=w_clk_cpu, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(22[6:15])
    
    wire n41467, n41516;
    wire [1:0]selected_1__N_340;
    
    wire w_clk_cpu_enable_547, n41456, n41458, n6, n24595;
    
    LUT4 i28976_2_lut_4_lut_4_lut (.A(n41426), .B(n41405), .C(n41467), 
         .D(n41424), .Z(n31536)) /* synthesis lut_function=(A (B)+!A (B ((D)+!C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(287[2] 289[5])
    defparam i28976_2_lut_4_lut_4_lut.init = 16'hcc8c;
    LUT4 equal_14_i3_2_lut_rep_429 (.A(selected[0]), .B(selected[1]), .Z(n41516)) /* synthesis lut_function=(A+(B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(253[7:20])
    defparam equal_14_i3_2_lut_rep_429.init = 16'heeee;
    LUT4 i28834_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(\selected_1__N_344[0] ), 
         .Z(selected_1__N_340[0])) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(253[7:20])
    defparam i28834_2_lut_3_lut.init = 16'h1010;
    LUT4 i37846_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(\selected_1__N_344[0] ), 
         .Z(selected_1__N_340[1])) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(253[7:20])
    defparam i37846_2_lut_3_lut.init = 16'h0101;
    FD1P3AX selected_i0 (.D(selected_1__N_340[0]), .SP(w_clk_cpu_enable_547), 
            .CK(w_clk_cpu), .Q(selected[0])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=1, LSE_RCOL=20, LSE_LLINE=451, LSE_RLINE=492 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(252[7] 275[5])
    defparam selected_i0.GSR = "ENABLED";
    LUT4 i29259_3_lut_rep_369_4_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_SEL_O[3]), 
         .D(LM32D_SEL_O[2]), .Z(n41456)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i29259_3_lut_rep_369_4_lut.init = 16'h4440;
    LUT4 i28838_2_lut_rep_363_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_WE_O), 
         .Z(w_clk_cpu_enable_303)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i28838_2_lut_rep_363_3_lut.init = 16'h4040;
    LUT4 i37901_2_lut_3_lut_4_lut (.A(selected[0]), .B(selected[1]), .C(n92[0]), 
         .D(LM32D_WE_O), .Z(n39983)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i37901_2_lut_3_lut_4_lut.init = 16'hbfff;
    LUT4 WBS_ADR_I_31__I_0_i12_4_lut_4_lut (.A(\LM32I_ADR_O[11] ), .B(\LM32D_ADR_O[11] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[11] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i12_4_lut_4_lut.init = 16'h0ca0;
    LUT4 i1_2_lut_rep_305_3_lut_4_lut_4_lut (.A(LM32D_SEL_O[2]), .B(selected[0]), 
         .C(selected[1]), .D(n25515), .Z(n41392)) /* synthesis lut_function=(A (B (C (D))+!B !(C+!(D)))+!A (B (C (D))+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(288[2] 289[4])
    defparam i1_2_lut_rep_305_3_lut_4_lut_4_lut.init = 16'hd300;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(LM32D_SEL_O[2]), .B(selected[0]), 
         .C(selected[1]), .D(n38761), .Z(PIO_OUT_15__N_3318)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(288[2] 289[4])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h2c00;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_432 (.A(LM32D_SEL_O[2]), .B(selected[0]), 
         .C(selected[1]), .D(n41344), .Z(n22230)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C (D)))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(288[2] 289[4])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_432.init = 16'h2c00;
    LUT4 WBS_ADR_I_31__I_0_i6_4_lut_4_lut (.A(\LM32I_ADR_O[5] ), .B(\LM32D_ADR_O[5] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[5] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i6_4_lut_4_lut.init = 16'h0ca0;
    LUT4 WBS_ADR_I_31__I_0_i9_4_lut_4_lut (.A(\LM32I_ADR_O[8] ), .B(\LM32D_ADR_O[8] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[8] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i9_4_lut_4_lut.init = 16'h0ca0;
    LUT4 WBS_ADR_I_31__I_0_i13_4_lut_4_lut (.A(\LM32I_ADR_O[12] ), .B(\LM32D_ADR_O[12] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[12] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i13_4_lut_4_lut.init = 16'h0ca0;
    LUT4 i23487_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(w_clk_cpu_enable_900), 
         .Z(n26128)) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i23487_2_lut_3_lut.init = 16'hb0b0;
    LUT4 WBS_ADR_I_31__I_0_i18_4_lut_4_lut (.A(\LM32I_ADR_O[17] ), .B(\LM32D_ADR_O[17] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[17] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i18_4_lut_4_lut.init = 16'h0ca0;
    LUT4 i28836_2_lut_rep_371_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_SEL_O[0]), 
         .Z(n41458)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i28836_2_lut_rep_371_3_lut.init = 16'h4040;
    LUT4 WBS_ADR_I_31__I_0_i17_4_lut_4_lut (.A(\LM32I_ADR_O[16] ), .B(\LM32D_ADR_O[16] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[16] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i17_4_lut_4_lut.init = 16'h0ca0;
    LUT4 WBS_ADR_I_31__I_0_i19_4_lut_4_lut (.A(\LM32I_ADR_O[18] ), .B(\LM32D_ADR_O[18] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[18] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i19_4_lut_4_lut.init = 16'h0ca0;
    LUT4 WBS_ADR_I_31__I_0_i16_4_lut_4_lut (.A(\LM32I_ADR_O[15] ), .B(\LM32D_ADR_O[15] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[15] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i16_4_lut_4_lut.init = 16'h0ca0;
    LUT4 WBS_ADR_I_31__I_0_i15_4_lut_4_lut (.A(\LM32I_ADR_O[14] ), .B(\LM32D_ADR_O[14] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[14] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i15_4_lut_4_lut.init = 16'h0ca0;
    LUT4 i29043_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(\LM32D_DAT_O[24] ), 
         .Z(\SHAREDBUS_DAT_I[24] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i29043_2_lut_3_lut.init = 16'h4040;
    LUT4 i28992_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(\LM32D_DAT_O[25] ), 
         .Z(\SHAREDBUS_DAT_I[25] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i28992_2_lut_3_lut.init = 16'h4040;
    LUT4 i28852_2_lut_3_lut_4_lut_3_lut (.A(selected[0]), .B(selected[1]), 
         .C(LM32D_SEL_O[1]), .Z(\SHAREDBUS_SEL_I[1] )) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i28852_2_lut_3_lut_4_lut_3_lut.init = 16'h6262;
    LUT4 i37871_2_lut_rep_339_3_lut_3_lut_4_lut_3_lut (.A(selected[0]), .B(selected[1]), 
         .C(LM32D_SEL_O[0]), .Z(n41426)) /* synthesis lut_function=(A (B)+!A !(B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i37871_2_lut_rep_339_3_lut_3_lut_4_lut_3_lut.init = 16'h9d9d;
    LUT4 i28839_2_lut_rep_342_3_lut_4_lut_3_lut (.A(selected[0]), .B(selected[1]), 
         .C(LM32D_SEL_O[2]), .Z(n41429)) /* synthesis lut_function=(!(A (B)+!A !(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i28839_2_lut_rep_342_3_lut_4_lut_3_lut.init = 16'h6262;
    LUT4 WBS_ADR_I_31__I_0_i20_4_lut_4_lut (.A(\LM32I_ADR_O[19] ), .B(\LM32D_ADR_O[19] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[19] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i20_4_lut_4_lut.init = 16'h0ca0;
    LUT4 WBS_ADR_I_31__I_0_i8_4_lut_4_lut (.A(\LM32I_ADR_O[7] ), .B(\LM32D_ADR_O[7] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[7] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i8_4_lut_4_lut.init = 16'h0ca0;
    LUT4 WBS_ADR_I_31__I_0_i11_4_lut_4_lut (.A(\LM32I_ADR_O[10] ), .B(\LM32D_ADR_O[10] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[10] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i11_4_lut_4_lut.init = 16'h0ca0;
    LUT4 WBS_ADR_I_31__I_0_i10_4_lut_4_lut (.A(\LM32I_ADR_O[9] ), .B(\LM32D_ADR_O[9] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[9] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i10_4_lut_4_lut.init = 16'h0ca0;
    LUT4 WBS_ADR_I_31__I_0_i7_4_lut_4_lut (.A(\LM32I_ADR_O[6] ), .B(\LM32D_ADR_O[6] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[6] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i7_4_lut_4_lut.init = 16'h0ca0;
    LUT4 i2_2_lut_3_lut_4_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_SEL_O[3]), 
         .D(LM32D_SEL_O[1]), .Z(n6)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 WBS_ADR_I_31__I_0_i5_4_lut_4_lut (.A(\LM32I_ADR_O[4] ), .B(\LM32D_ADR_O[4] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[4] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i5_4_lut_4_lut.init = 16'h0ca0;
    LUT4 WBS_ADR_I_31__I_0_i32_4_lut_rep_355_4_lut (.A(\LM32I_ADR_O[31] ), 
         .B(\LM32D_ADR_O[31] ), .C(selected[0]), .D(selected[1]), .Z(n41442)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i32_4_lut_rep_355_4_lut.init = 16'h0ca0;
    LUT4 i38066_2_lut_rep_336_3_lut_3_lut_4_lut_3_lut (.A(selected[0]), .B(selected[1]), 
         .C(LM32D_SEL_O[3]), .Z(n41423)) /* synthesis lut_function=(A (B)+!A !(B (C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i38066_2_lut_rep_336_3_lut_3_lut_4_lut_3_lut.init = 16'h9d9d;
    LUT4 WBS_ADR_I_31__I_0_i14_4_lut_rep_348_4_lut (.A(\LM32I_ADR_O[13] ), 
         .B(\LM32D_ADR_O[13] ), .C(selected[0]), .D(selected[1]), .Z(n41435)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i14_4_lut_rep_348_4_lut.init = 16'h0ca0;
    LUT4 WBS_ADR_I_31__I_0_i23_4_lut_4_lut (.A(\LM32I_ADR_O[22] ), .B(\LM32D_ADR_O[22] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[22] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i23_4_lut_4_lut.init = 16'h0ca0;
    LUT4 WBS_ADR_I_31__I_0_i27_4_lut_4_lut (.A(\LM32I_ADR_O[26] ), .B(\LM32D_ADR_O[26] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[26] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i27_4_lut_4_lut.init = 16'h0ca0;
    LUT4 WBS_ADR_I_31__I_0_i26_4_lut_4_lut (.A(\LM32I_ADR_O[25] ), .B(\LM32D_ADR_O[25] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[25] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i26_4_lut_4_lut.init = 16'h0ca0;
    LUT4 WBS_ADR_I_31__I_0_i25_4_lut_4_lut (.A(\LM32I_ADR_O[24] ), .B(\LM32D_ADR_O[24] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[24] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i25_4_lut_4_lut.init = 16'h0ca0;
    LUT4 WBS_ADR_I_31__I_0_i28_4_lut_4_lut (.A(\LM32I_ADR_O[27] ), .B(\LM32D_ADR_O[27] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[27] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i28_4_lut_4_lut.init = 16'h0ca0;
    LUT4 WBS_ADR_I_31__I_0_i29_4_lut_4_lut (.A(\LM32I_ADR_O[28] ), .B(\LM32D_ADR_O[28] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[28] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i29_4_lut_4_lut.init = 16'h0ca0;
    LUT4 i28984_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(\LM32D_DAT_O[26] ), 
         .Z(\SHAREDBUS_DAT_I[26] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i28984_2_lut_3_lut.init = 16'h4040;
    LUT4 i28902_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(\LM32D_DAT_O[28] ), 
         .Z(\SHAREDBUS_DAT_I[28] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i28902_2_lut_3_lut.init = 16'h4040;
    LUT4 WBS_ADR_I_31__I_0_i30_4_lut_4_lut (.A(\LM32I_ADR_O[29] ), .B(\LM32D_ADR_O[29] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[29] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i30_4_lut_4_lut.init = 16'h0ca0;
    LUT4 i28894_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(\LM32D_DAT_O[29] ), 
         .Z(\SHAREDBUS_DAT_I[29] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i28894_2_lut_3_lut.init = 16'h4040;
    LUT4 i28885_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(\LM32D_DAT_O[30] ), 
         .Z(\SHAREDBUS_DAT_I[30] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i28885_2_lut_3_lut.init = 16'h4040;
    LUT4 i28884_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(\LM32D_DAT_O[31] ), 
         .Z(\SHAREDBUS_DAT_I[31] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i28884_2_lut_3_lut.init = 16'h4040;
    LUT4 i29173_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(\LM32D_DAT_O[18] ), 
         .Z(\SHAREDBUS_DAT_I[18] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i29173_2_lut_3_lut.init = 16'h4040;
    LUT4 i29149_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(\LM32D_DAT_O[19] ), 
         .Z(\SHAREDBUS_DAT_I[19] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i29149_2_lut_3_lut.init = 16'h4040;
    LUT4 WBS_ADR_I_31__I_0_i24_4_lut_4_lut (.A(\LM32I_ADR_O[23] ), .B(\LM32D_ADR_O[23] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[23] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i24_4_lut_4_lut.init = 16'h0ca0;
    LUT4 WBS_ADR_I_31__I_0_i31_4_lut_4_lut (.A(\LM32I_ADR_O[30] ), .B(\LM32D_ADR_O[30] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[30] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i31_4_lut_4_lut.init = 16'h0ca0;
    LUT4 i29078_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(\LM32D_DAT_O[20] ), 
         .Z(\SHAREDBUS_DAT_I[20] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i29078_2_lut_3_lut.init = 16'h4040;
    LUT4 WBS_ADR_I_31__I_0_i22_4_lut_4_lut (.A(\LM32I_ADR_O[21] ), .B(\LM32D_ADR_O[21] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[21] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i22_4_lut_4_lut.init = 16'h0ca0;
    LUT4 WBS_ADR_I_31__I_0_i3_4_lut_4_lut (.A(\LM32I_ADR_O[2] ), .B(\LM32D_ADR_O[2] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[2] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i3_4_lut_4_lut.init = 16'h0ca0;
    LUT4 i29075_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(\LM32D_DAT_O[21] ), 
         .Z(\SHAREDBUS_DAT_I[21] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i29075_2_lut_3_lut.init = 16'h4040;
    LUT4 WBS_ADR_I_31__I_0_i4_4_lut_4_lut (.A(\LM32I_ADR_O[3] ), .B(\LM32D_ADR_O[3] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[3] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i4_4_lut_4_lut.init = 16'h0ca0;
    LUT4 i29063_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(\LM32D_DAT_O[22] ), 
         .Z(\SHAREDBUS_DAT_I[22] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i29063_2_lut_3_lut.init = 16'h4040;
    LUT4 i29044_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(\LM32D_DAT_O[23] ), 
         .Z(\SHAREDBUS_DAT_I[23] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i29044_2_lut_3_lut.init = 16'h4040;
    LUT4 i28950_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(\LM32D_DAT_O[27] ), 
         .Z(\SHAREDBUS_DAT_I[27] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i28950_2_lut_3_lut.init = 16'h4040;
    LUT4 WBS_ADR_I_31__I_0_i21_4_lut_4_lut (.A(\LM32I_ADR_O[20] ), .B(\LM32D_ADR_O[20] ), 
         .C(selected[0]), .D(selected[1]), .Z(\SHAREDBUS_ADR_I[20] )) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(279[2] 281[5])
    defparam WBS_ADR_I_31__I_0_i21_4_lut_4_lut.init = 16'h0ca0;
    LUT4 mux_18_i1_4_lut_4_lut (.A(LM32I_CYC_O), .B(LM32D_CYC_O), .C(selected[0]), 
         .D(selected[1]), .Z(n92[0])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(307[2] 309[5])
    defparam mux_18_i1_4_lut_4_lut.init = 16'h0ca0;
    LUT4 mux_19_i1_4_lut_4_lut (.A(\selected_1__N_344[0] ), .B(LM32D_STB_O), 
         .C(selected[0]), .D(selected[1]), .Z(n93[0])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B ((D)+!C))+!A ((C+!(D))+!B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(311[2] 313[5])
    defparam mux_19_i1_4_lut_4_lut.init = 16'h0ca0;
    LUT4 i2_3_lut_4_lut (.A(n41479), .B(n41456), .C(n41458), .D(n41467), 
         .Z(n38998)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(287[2] 289[5])
    defparam i2_3_lut_4_lut.init = 16'hffef;
    LUT4 i2_3_lut_rep_306_3_lut_4_lut (.A(n41479), .B(n41456), .C(n41467), 
         .D(n41426), .Z(n41393)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(287[2] 289[5])
    defparam i2_3_lut_rep_306_3_lut_4_lut.init = 16'hffef;
    FD1P3AX selected_i1 (.D(selected_1__N_340[1]), .SP(w_clk_cpu_enable_547), 
            .CK(w_clk_cpu), .Q(selected[1])) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=1, LSE_RCOL=20, LSE_LLINE=451, LSE_RLINE=492 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(252[7] 275[5])
    defparam selected_i1.GSR = "ENABLED";
    LUT4 i28882_2_lut_rep_380_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_SEL_O[1]), 
         .Z(n41467)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i28882_2_lut_rep_380_3_lut.init = 16'h4040;
    LUT4 mux_8_i4_3_lut_4_lut (.A(n41469), .B(n41479), .C(\SHAREDBUS_DAT_I[19] ), 
         .D(\data[19] ), .Z(n87[3])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(287[2] 289[5])
    defparam mux_8_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i37896_2_lut_rep_276_2_lut_3_lut_4_lut (.A(n41469), .B(n41479), 
         .C(n41390), .D(n25515), .Z(n41363)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+(D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(287[2] 289[5])
    defparam i37896_2_lut_rep_276_2_lut_3_lut_4_lut.init = 16'h0e0f;
    LUT4 mux_8_i1_3_lut_4_lut (.A(n41469), .B(n41479), .C(\SHAREDBUS_DAT_I[16] ), 
         .D(\data[16] ), .Z(n87[0])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(287[2] 289[5])
    defparam mux_8_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_8_i2_3_lut_4_lut (.A(n41469), .B(n41479), .C(\SHAREDBUS_DAT_I[17] ), 
         .D(\data[17] ), .Z(n87[1])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(287[2] 289[5])
    defparam mux_8_i2_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_8_i8_3_lut_4_lut (.A(n41469), .B(n41479), .C(\SHAREDBUS_DAT_I[23] ), 
         .D(\data[23] ), .Z(n87[7])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(287[2] 289[5])
    defparam mux_8_i8_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_8_i3_3_lut_4_lut (.A(n41469), .B(n41479), .C(\SHAREDBUS_DAT_I[18] ), 
         .D(\data[18] ), .Z(n87[2])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(287[2] 289[5])
    defparam mux_8_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_8_i7_3_lut_4_lut (.A(n41469), .B(n41479), .C(\SHAREDBUS_DAT_I[22] ), 
         .D(\data[22] ), .Z(n87[6])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(287[2] 289[5])
    defparam mux_8_i7_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_8_i5_3_lut_4_lut (.A(n41469), .B(n41479), .C(\SHAREDBUS_DAT_I[20] ), 
         .D(\data[20] ), .Z(n87[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(287[2] 289[5])
    defparam mux_8_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_8_i6_3_lut_4_lut (.A(n41469), .B(n41479), .C(\SHAREDBUS_DAT_I[21] ), 
         .D(\data[21] ), .Z(n87[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(287[2] 289[5])
    defparam mux_8_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i2_4_lut_rep_303_4_lut (.A(n41426), .B(n41490), .C(n24709), .D(\SHAREDBUS_SEL_I[1] ), 
         .Z(n41390)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(287[2] 289[5])
    defparam i2_4_lut_rep_303_4_lut.init = 16'h0020;
    LUT4 i37907_4_lut_rep_318 (.A(n41479), .B(n41458), .C(n6), .D(LM32D_SEL_O[2]), 
         .Z(n41405)) /* synthesis lut_function=(!(A+(B (C (D))))) */ ;
    defparam i37907_4_lut_rep_318.init = 16'h1555;
    LUT4 i37934_2_lut_rep_325_2_lut_3_lut_2_lut (.A(selected[0]), .B(selected[1]), 
         .Z(n41412)) /* synthesis lut_function=(!(A+!(B))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i37934_2_lut_rep_325_2_lut_3_lut_2_lut.init = 16'h4444;
    LUT4 i28861_2_lut_rep_368_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_SEL_O[3]), 
         .Z(n41455)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i28861_2_lut_rep_368_3_lut.init = 16'h4040;
    LUT4 i29299_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(\LM32D_DAT_O[17] ), 
         .Z(\SHAREDBUS_DAT_I[17] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i29299_2_lut_3_lut.init = 16'h4040;
    LUT4 \genblk5.tmp_ack_o_d_I_0_3_lut_rep_334_4_lut  (.A(LM32D_WE_O), .B(n41490), 
         .C(tmp_ack_o), .D(\genblk5.tmp_ack_o_d ), .Z(n41421)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(292[2] 293[4])
    defparam \genblk5.tmp_ack_o_d_I_0_3_lut_rep_334_4_lut .init = 16'hfd20;
    LUT4 i2_3_lut_4_lut_adj_433 (.A(LM32D_WE_O), .B(n41490), .C(n42723), 
         .D(n25664), .Z(n36688)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(292[2] 293[4])
    defparam i2_3_lut_4_lut_adj_433.init = 16'h0020;
    LUT4 i21682_2_lut_3_lut_3_lut_4_lut_4_lut (.A(n41479), .B(n41429), .C(n25515), 
         .D(n41458), .Z(n24342)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C (D))))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(316[22:38])
    defparam i21682_2_lut_3_lut_3_lut_4_lut_4_lut.init = 16'h3020;
    LUT4 n20799_bdd_2_lut_3_lut_4_lut_4_lut (.A(n41479), .B(n25515), .C(n41429), 
         .D(n41458), .Z(n36822)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(316[22:38])
    defparam n20799_bdd_2_lut_3_lut_4_lut_4_lut.init = 16'hfffb;
    LUT4 i2_3_lut_4_lut_4_lut (.A(n41479), .B(n41456), .C(\SHAREDBUS_SEL_I[1] ), 
         .D(n41458), .Z(n37005)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(316[22:38])
    defparam i2_3_lut_4_lut_4_lut.init = 16'h0010;
    LUT4 i29366_2_lut_3_lut (.A(selected[0]), .B(selected[1]), .C(\LM32D_DAT_O[16] ), 
         .Z(\SHAREDBUS_DAT_I[16] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i29366_2_lut_3_lut.init = 16'h4040;
    LUT4 i28864_2_lut_rep_382_3_lut (.A(selected[0]), .B(selected[1]), .C(LM32D_SEL_O[2]), 
         .Z(n41469)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i28864_2_lut_rep_382_3_lut.init = 16'h4040;
    LUT4 i1_3_lut_4_lut (.A(\selected_1__N_344[0] ), .B(n41516), .C(LM32D_STB_O), 
         .D(n24595), .Z(w_clk_cpu_enable_547)) /* synthesis lut_function=(A ((D)+!B)+!A (B (D)+!B (C))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hfe32;
    LUT4 i21972_4_lut_4_lut (.A(n41479), .B(n41352), .C(n41490), .D(n76[0]), 
         .Z(n24595)) /* synthesis lut_function=(A (B+(D))+!A !(B (C)+!B (C+!(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(316[22:38])
    defparam i21972_4_lut_4_lut.init = 16'haf8c;
    LUT4 i2_3_lut_4_lut_4_lut_adj_434 (.A(LM32D_SEL_O[2]), .B(n41490), .C(n39016), 
         .D(LM32D_SEL_O[3]), .Z(n39018)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(288[2] 289[4])
    defparam i2_3_lut_4_lut_4_lut_adj_434.init = 16'hfeff;
    LUT4 i26064_4_lut (.A(n21531), .B(\sramsram_data_in[3] ), .C(n7), 
         .D(n28684), .Z(\tmp_dat_o_nxt_31__N_3207[19] )) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i26064_4_lut.init = 16'hca0a;
    LUT4 selected_1__I_0_i3_2_lut_rep_403 (.A(selected[0]), .B(selected[1]), 
         .Z(n41490)) /* synthesis lut_function=(A+!(B)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam selected_1__I_0_i3_2_lut_rep_403.init = 16'hbbbb;
    LUT4 i37972_2_lut_rep_392 (.A(selected[0]), .B(selected[1]), .Z(n41479)) /* synthesis lut_function=(!((B)+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(316[22:38])
    defparam i37972_2_lut_rep_392.init = 16'h2222;
    LUT4 i2_3_lut_3_lut_4_lut (.A(selected[0]), .B(selected[1]), .C(n38871), 
         .D(LM32I_CYC_O), .Z(bus_error_f_N_1764)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(316[22:38])
    defparam i2_3_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i29185_2_lut_3_lut_3_lut_4_lut_3_lut (.A(selected[0]), .B(selected[1]), 
         .C(\LM32D_ADR_O[0] ), .Z(\SHAREDBUS_ADR_I[0] )) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/mico_cpu/soc/mico_cpu.v(321[22:38])
    defparam i29185_2_lut_3_lut_3_lut_4_lut_3_lut.init = 16'h4040;
    
endmodule
//
// Verilog Description of module lm32_top
//

module lm32_top (GND_net, n41435, n7, n7_adj_64, n7_adj_65, n7_adj_66, 
            n7_adj_67, n7_adj_68, n7_adj_69, n7_adj_70, n7_adj_71, 
            n7_adj_72, n7_adj_73, n7_adj_74, n7_adj_75, n7_adj_76, 
            n7_adj_77, n7_adj_78, n7_adj_79, n7_adj_80, n7_adj_81, 
            n7_adj_82, n7_adj_83, n7_adj_84, n7_adj_85, n7_adj_86, 
            n7_adj_87, n7_adj_88, n7_adj_89, n7_adj_90, n7_adj_91, 
            n7_adj_92, n7_adj_93, n7_adj_94, LM32DEBUG_ACK_O, w_result, 
            w_clk_cpu, data_bus_error_exception_N_1225, n42726, read_idx_0_d, 
            n23059, n23091, n23058, n23090, n23067, n23099, LM32D_CYC_O, 
            n23068, n23100, LM32I_CYC_O, n42734, n42738, read_idx_1_d, 
            n23069, n23101, n42732, n23070, n23102, n23071, n23103, 
            n23072, n23104, \counter[2] , n41470, write_idx_w, n23185, 
            n23186, n23073, n23105, n23074, n23106, n23075, n23107, 
            n23076, n23108, n22885, wb_load_complete_N_2129, reg_data_1, 
            n23056, n23088, n23057, n23089, n22999, n22877, n22874, 
            n23053, n23085, n23054, n23086, n23060, n23092, n23061, 
            n23093, n23062, n23094, n23063, n23095, n23064, n23096, 
            n23065, n23097, n23066, n23098, n23052, n23084, n23055, 
            n23087, n23077, n23109, n23078, n23110, n23079, n23111, 
            n23080, n23112, n23081, n23113, n23082, n23114, n23083, 
            n23115, i_cyc_o_N_1759, LM32D_WE_O, LM32D_DAT_O, SHAREDBUS_DAT_O, 
            LM32D_ADR_O, LM32D_SEL_O, LM32D_STB_O, \LM32I_ADR_O[2] , 
            \selected_1__N_344[0] , \LM32I_ADR_O[31] , bus_error_f_N_1764, 
            \LM32I_ADR_O[30] , \LM32I_ADR_O[29] , \LM32I_ADR_O[28] , \LM32I_ADR_O[27] , 
            \LM32I_ADR_O[26] , \LM32I_ADR_O[25] , \LM32I_ADR_O[24] , \LM32I_ADR_O[23] , 
            \LM32I_ADR_O[22] , \LM32I_ADR_O[21] , \LM32I_ADR_O[20] , \LM32I_ADR_O[19] , 
            \LM32I_ADR_O[18] , \LM32I_ADR_O[17] , \LM32I_ADR_O[16] , \LM32I_ADR_O[15] , 
            \LM32I_ADR_O[14] , \LM32I_ADR_O[13] , \LM32I_ADR_O[12] , \LM32I_ADR_O[11] , 
            \LM32I_ADR_O[10] , \LM32I_ADR_O[9] , \LM32I_ADR_O[8] , \LM32I_ADR_O[7] , 
            \LM32I_ADR_O[6] , \LM32I_ADR_O[5] , \LM32I_ADR_O[4] , \LM32I_ADR_O[3] , 
            n41479, n38871, \data[31] , n87, \SHAREDBUS_SEL_I[1] , 
            n41490, \data[21] , \data[19] , w_clk_cpu_enable_303, \data[30] , 
            n41426, \data[29] , \data[28] , n93, n92, n41422, n35, 
            \data[27] , \data[26] , \data[25] , \data[18] , \data[24] , 
            \data[23] , \data[17] , \data[16] , n96, \data[22] , \data[20] , 
            \SHAREDBUS_ADR_I[10] , \SHAREDBUS_ADR_I[9] , \SHAREDBUS_ADR_I[8] , 
            \SHAREDBUS_ADR_I[7] , \SHAREDBUS_ADR_I[6] , \SHAREDBUS_ADR_I[5] , 
            \SHAREDBUS_ADR_I[4] , \SHAREDBUS_ADR_I[3] , \SHAREDBUS_ADR_I[2] , 
            VCC_net, counter_2__N_178) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    input n41435;
    output n7;
    output n7_adj_64;
    output n7_adj_65;
    output n7_adj_66;
    output n7_adj_67;
    output n7_adj_68;
    output n7_adj_69;
    output n7_adj_70;
    output n7_adj_71;
    output n7_adj_72;
    output n7_adj_73;
    output n7_adj_74;
    output n7_adj_75;
    output n7_adj_76;
    output n7_adj_77;
    output n7_adj_78;
    output n7_adj_79;
    output n7_adj_80;
    output n7_adj_81;
    output n7_adj_82;
    output n7_adj_83;
    output n7_adj_84;
    output n7_adj_85;
    output n7_adj_86;
    output n7_adj_87;
    output n7_adj_88;
    output n7_adj_89;
    output n7_adj_90;
    output n7_adj_91;
    output n7_adj_92;
    output n7_adj_93;
    output n7_adj_94;
    output LM32DEBUG_ACK_O;
    output [31:0]w_result;
    input w_clk_cpu;
    input data_bus_error_exception_N_1225;
    input n42726;
    output [4:0]read_idx_0_d;
    input n23059;
    input n23091;
    input n23058;
    input n23090;
    input n23067;
    input n23099;
    output LM32D_CYC_O;
    input n23068;
    input n23100;
    output LM32I_CYC_O;
    output n42734;
    output n42738;
    output [4:0]read_idx_1_d;
    input n23069;
    input n23101;
    output n42732;
    input n23070;
    input n23102;
    input n23071;
    input n23103;
    input n23072;
    input n23104;
    input \counter[2] ;
    output n41470;
    output [4:0]write_idx_w;
    output n23185;
    output n23186;
    input n23073;
    input n23105;
    input n23074;
    input n23106;
    input n23075;
    input n23107;
    input n23076;
    input n23108;
    input n22885;
    input wb_load_complete_N_2129;
    input [31:0]reg_data_1;
    input n23056;
    input n23088;
    input n23057;
    input n23089;
    input n22999;
    output n22877;
    output n22874;
    input n23053;
    input n23085;
    input n23054;
    input n23086;
    input n23060;
    input n23092;
    input n23061;
    input n23093;
    input n23062;
    input n23094;
    input n23063;
    input n23095;
    input n23064;
    input n23096;
    input n23065;
    input n23097;
    input n23066;
    input n23098;
    input n23052;
    input n23084;
    input n23055;
    input n23087;
    input n23077;
    input n23109;
    input n23078;
    input n23110;
    input n23079;
    input n23111;
    input n23080;
    input n23112;
    input n23081;
    input n23113;
    input n23082;
    input n23114;
    input n23083;
    input n23115;
    input i_cyc_o_N_1759;
    output LM32D_WE_O;
    output [31:0]LM32D_DAT_O;
    input [31:0]SHAREDBUS_DAT_O;
    output [31:0]LM32D_ADR_O;
    output [3:0]LM32D_SEL_O;
    output LM32D_STB_O;
    output \LM32I_ADR_O[2] ;
    output \selected_1__N_344[0] ;
    output \LM32I_ADR_O[31] ;
    input bus_error_f_N_1764;
    output \LM32I_ADR_O[30] ;
    output \LM32I_ADR_O[29] ;
    output \LM32I_ADR_O[28] ;
    output \LM32I_ADR_O[27] ;
    output \LM32I_ADR_O[26] ;
    output \LM32I_ADR_O[25] ;
    output \LM32I_ADR_O[24] ;
    output \LM32I_ADR_O[23] ;
    output \LM32I_ADR_O[22] ;
    output \LM32I_ADR_O[21] ;
    output \LM32I_ADR_O[20] ;
    output \LM32I_ADR_O[19] ;
    output \LM32I_ADR_O[18] ;
    output \LM32I_ADR_O[17] ;
    output \LM32I_ADR_O[16] ;
    output \LM32I_ADR_O[15] ;
    output \LM32I_ADR_O[14] ;
    output \LM32I_ADR_O[13] ;
    output \LM32I_ADR_O[12] ;
    output \LM32I_ADR_O[11] ;
    output \LM32I_ADR_O[10] ;
    output \LM32I_ADR_O[9] ;
    output \LM32I_ADR_O[8] ;
    output \LM32I_ADR_O[7] ;
    output \LM32I_ADR_O[6] ;
    output \LM32I_ADR_O[5] ;
    output \LM32I_ADR_O[4] ;
    output \LM32I_ADR_O[3] ;
    input n41479;
    input n38871;
    output \data[31] ;
    input [7:0]n87;
    input \SHAREDBUS_SEL_I[1] ;
    input n41490;
    output \data[21] ;
    output \data[19] ;
    input w_clk_cpu_enable_303;
    output \data[30] ;
    input n41426;
    output \data[29] ;
    output \data[28] ;
    input [0:0]n93;
    input [0:0]n92;
    output n41422;
    input n35;
    output \data[27] ;
    output \data[26] ;
    output \data[25] ;
    output \data[18] ;
    output \data[24] ;
    output \data[23] ;
    output \data[17] ;
    output \data[16] ;
    input [7:0]n96;
    output \data[22] ;
    output \data[20] ;
    input \SHAREDBUS_ADR_I[10] ;
    input \SHAREDBUS_ADR_I[9] ;
    input \SHAREDBUS_ADR_I[8] ;
    input \SHAREDBUS_ADR_I[7] ;
    input \SHAREDBUS_ADR_I[6] ;
    input \SHAREDBUS_ADR_I[5] ;
    input \SHAREDBUS_ADR_I[4] ;
    input \SHAREDBUS_ADR_I[3] ;
    input \SHAREDBUS_ADR_I[2] ;
    input VCC_net;
    input counter_2__N_178;
    
    wire jtag_update_N_2932 /* synthesis is_inv_clock=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(203[14:23])
    wire jtag_update /* synthesis is_clock=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(254[6:17])
    wire w_clk_cpu /* synthesis SET_AS_NETWORK=w_clk_cpu, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(22[6:15])
    wire [7:0]jtag_reg_d;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(248[23:33])
    wire [7:0]jtag_reg_q;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(252[12:22])
    wire [2:0]jtag_reg_addr_d;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(255[12:27])
    wire [2:0]jtag_reg_addr_q;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(256[12:27])
    wire [31:0]ROM_DAT_O;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(392[26:35])
    
    wire ROM_ACK_O;
    
    INV i39325 (.A(jtag_update), .Z(jtag_update_N_2932));
    jtag_cores jtag_cores (.reg_d({jtag_reg_d}), .reg_addr_d({GND_net, jtag_reg_addr_d[1:0]}), 
            .reg_update(jtag_update), .reg_q({jtag_reg_q}), .reg_addr_q({jtag_reg_addr_q})) /* synthesis LSE_LINE_FILE_ID=8, LSE_LCOL=2, LSE_RCOL=36, LSE_LLINE=519, LSE_RLINE=560, syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(418[12] 432[6])
    LUT4 i1_2_lut_2_lut (.A(n41435), .B(ROM_DAT_O[5]), .Z(n7)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_401 (.A(n41435), .B(ROM_DAT_O[6]), .Z(n7_adj_64)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_401.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_402 (.A(n41435), .B(ROM_DAT_O[7]), .Z(n7_adj_65)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_402.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_403 (.A(n41435), .B(ROM_DAT_O[8]), .Z(n7_adj_66)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_403.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_404 (.A(n41435), .B(ROM_DAT_O[9]), .Z(n7_adj_67)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_404.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_405 (.A(n41435), .B(ROM_DAT_O[11]), .Z(n7_adj_68)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_405.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_406 (.A(n41435), .B(ROM_DAT_O[12]), .Z(n7_adj_69)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_406.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_407 (.A(n41435), .B(ROM_DAT_O[13]), .Z(n7_adj_70)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_407.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_408 (.A(n41435), .B(ROM_DAT_O[14]), .Z(n7_adj_71)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_408.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_409 (.A(n41435), .B(ROM_DAT_O[15]), .Z(n7_adj_72)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_409.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_410 (.A(n41435), .B(ROM_DAT_O[16]), .Z(n7_adj_73)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_410.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_411 (.A(n41435), .B(ROM_DAT_O[17]), .Z(n7_adj_74)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_411.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_412 (.A(n41435), .B(ROM_DAT_O[18]), .Z(n7_adj_75)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_412.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_413 (.A(n41435), .B(ROM_DAT_O[19]), .Z(n7_adj_76)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_413.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_414 (.A(n41435), .B(ROM_DAT_O[20]), .Z(n7_adj_77)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_414.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_415 (.A(n41435), .B(ROM_DAT_O[21]), .Z(n7_adj_78)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_415.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_416 (.A(n41435), .B(ROM_DAT_O[22]), .Z(n7_adj_79)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_416.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_417 (.A(n41435), .B(ROM_DAT_O[23]), .Z(n7_adj_80)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_417.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_418 (.A(n41435), .B(ROM_DAT_O[24]), .Z(n7_adj_81)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_418.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_419 (.A(n41435), .B(ROM_DAT_O[25]), .Z(n7_adj_82)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_419.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_420 (.A(n41435), .B(ROM_DAT_O[26]), .Z(n7_adj_83)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_420.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_421 (.A(n41435), .B(ROM_DAT_O[27]), .Z(n7_adj_84)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_421.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_422 (.A(n41435), .B(ROM_DAT_O[29]), .Z(n7_adj_85)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_422.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_423 (.A(n41435), .B(ROM_DAT_O[30]), .Z(n7_adj_86)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_423.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_424 (.A(n41435), .B(ROM_DAT_O[31]), .Z(n7_adj_87)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_424.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_425 (.A(n41435), .B(ROM_DAT_O[28]), .Z(n7_adj_88)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_425.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_426 (.A(n41435), .B(ROM_DAT_O[10]), .Z(n7_adj_89)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_426.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_427 (.A(n41435), .B(ROM_DAT_O[4]), .Z(n7_adj_90)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_427.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_428 (.A(n41435), .B(ROM_DAT_O[1]), .Z(n7_adj_91)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_428.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_429 (.A(n41435), .B(ROM_DAT_O[0]), .Z(n7_adj_92)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_429.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_430 (.A(n41435), .B(ROM_DAT_O[2]), .Z(n7_adj_93)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_430.init = 16'h4444;
    LUT4 i1_2_lut_2_lut_adj_431 (.A(n41435), .B(ROM_DAT_O[3]), .Z(n7_adj_94)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i1_2_lut_2_lut_adj_431.init = 16'h4444;
    LUT4 i28865_2_lut_2_lut (.A(n41435), .B(ROM_ACK_O), .Z(LM32DEBUG_ACK_O)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(403[45:61])
    defparam i28865_2_lut_2_lut.init = 16'h4444;
    lm32_cpu cpu (.w_result({w_result}), .w_clk_cpu(w_clk_cpu), .data_bus_error_exception_N_1225(data_bus_error_exception_N_1225), 
            .n42726(n42726), .read_idx_0_d({read_idx_0_d}), .n23059(n23059), 
            .n23091(n23091), .n23058(n23058), .n23090(n23090), .n23067(n23067), 
            .n23099(n23099), .LM32D_CYC_O(LM32D_CYC_O), .n23068(n23068), 
            .n23100(n23100), .LM32I_CYC_O(LM32I_CYC_O), .n42734(n42734), 
            .n42738(n42738), .read_idx_1_d({read_idx_1_d}), .n23069(n23069), 
            .n23101(n23101), .n42732(n42732), .n23070(n23070), .n23102(n23102), 
            .n23071(n23071), .n23103(n23103), .n23072(n23072), .n23104(n23104), 
            .\counter[2] (\counter[2] ), .n41470(n41470), .write_idx_w({write_idx_w}), 
            .n23185(n23185), .n23186(n23186), .n23073(n23073), .n23105(n23105), 
            .n23074(n23074), .n23106(n23106), .n23075(n23075), .n23107(n23107), 
            .n23076(n23076), .n23108(n23108), .n22885(n22885), .\jtag_reg_addr_d[0] (jtag_reg_addr_d[0]), 
            .\jtag_reg_addr_d[1] (jtag_reg_addr_d[1]), .wb_load_complete_N_2129(wb_load_complete_N_2129), 
            .GND_net(GND_net), .reg_data_1({reg_data_1}), .n23056(n23056), 
            .n23088(n23088), .n23057(n23057), .n23089(n23089), .n22999(n22999), 
            .n22877(n22877), .n22874(n22874), .n23053(n23053), .n23085(n23085), 
            .n23054(n23054), .n23086(n23086), .n23060(n23060), .n23092(n23092), 
            .n23061(n23061), .n23093(n23093), .n23062(n23062), .n23094(n23094), 
            .n23063(n23063), .n23095(n23095), .n23064(n23064), .n23096(n23096), 
            .n23065(n23065), .n23097(n23097), .n23066(n23066), .n23098(n23098), 
            .n23052(n23052), .n23084(n23084), .n23055(n23055), .n23087(n23087), 
            .n23077(n23077), .n23109(n23109), .n23078(n23078), .n23110(n23110), 
            .n23079(n23079), .n23111(n23111), .n23080(n23080), .n23112(n23112), 
            .n23081(n23081), .n23113(n23113), .n23082(n23082), .n23114(n23114), 
            .n23083(n23083), .n23115(n23115), .i_cyc_o_N_1759(i_cyc_o_N_1759), 
            .LM32D_WE_O(LM32D_WE_O), .LM32D_DAT_O({LM32D_DAT_O}), .SHAREDBUS_DAT_O({SHAREDBUS_DAT_O}), 
            .LM32D_ADR_O({LM32D_ADR_O}), .LM32D_SEL_O({LM32D_SEL_O}), .LM32D_STB_O(LM32D_STB_O), 
            .jtag_reg_d({jtag_reg_d}), .jtag_reg_q({jtag_reg_q}), .jtag_update_N_2932(jtag_update_N_2932), 
            .jtag_reg_addr_q({jtag_reg_addr_q}), .\LM32I_ADR_O[2] (\LM32I_ADR_O[2] ), 
            .\selected_1__N_344[0] (\selected_1__N_344[0] ), .\LM32I_ADR_O[31] (\LM32I_ADR_O[31] ), 
            .bus_error_f_N_1764(bus_error_f_N_1764), .\LM32I_ADR_O[30] (\LM32I_ADR_O[30] ), 
            .\LM32I_ADR_O[29] (\LM32I_ADR_O[29] ), .\LM32I_ADR_O[28] (\LM32I_ADR_O[28] ), 
            .\LM32I_ADR_O[27] (\LM32I_ADR_O[27] ), .\LM32I_ADR_O[26] (\LM32I_ADR_O[26] ), 
            .\LM32I_ADR_O[25] (\LM32I_ADR_O[25] ), .\LM32I_ADR_O[24] (\LM32I_ADR_O[24] ), 
            .\LM32I_ADR_O[23] (\LM32I_ADR_O[23] ), .\LM32I_ADR_O[22] (\LM32I_ADR_O[22] ), 
            .\LM32I_ADR_O[21] (\LM32I_ADR_O[21] ), .\LM32I_ADR_O[20] (\LM32I_ADR_O[20] ), 
            .\LM32I_ADR_O[19] (\LM32I_ADR_O[19] ), .\LM32I_ADR_O[18] (\LM32I_ADR_O[18] ), 
            .\LM32I_ADR_O[17] (\LM32I_ADR_O[17] ), .\LM32I_ADR_O[16] (\LM32I_ADR_O[16] ), 
            .\LM32I_ADR_O[15] (\LM32I_ADR_O[15] ), .\LM32I_ADR_O[14] (\LM32I_ADR_O[14] ), 
            .\LM32I_ADR_O[13] (\LM32I_ADR_O[13] ), .\LM32I_ADR_O[12] (\LM32I_ADR_O[12] ), 
            .\LM32I_ADR_O[11] (\LM32I_ADR_O[11] ), .\LM32I_ADR_O[10] (\LM32I_ADR_O[10] ), 
            .\LM32I_ADR_O[9] (\LM32I_ADR_O[9] ), .\LM32I_ADR_O[8] (\LM32I_ADR_O[8] ), 
            .\LM32I_ADR_O[7] (\LM32I_ADR_O[7] ), .\LM32I_ADR_O[6] (\LM32I_ADR_O[6] ), 
            .\LM32I_ADR_O[5] (\LM32I_ADR_O[5] ), .\LM32I_ADR_O[4] (\LM32I_ADR_O[4] ), 
            .\LM32I_ADR_O[3] (\LM32I_ADR_O[3] ), .n41479(n41479), .n38871(n38871)) /* synthesis syn_module_defined=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(283[10] 366[6])
    lm32_monitor ROM_DAT_O_31__I_13 (.data({\data[31] , Open_7, Open_8, 
            Open_9, Open_10, Open_11, Open_12, Open_13, Open_14, 
            Open_15, Open_16, Open_17, Open_18, Open_19, Open_20, 
            Open_21, Open_22, Open_23, Open_24, Open_25, Open_26, 
            Open_27, Open_28, Open_29, Open_30, Open_31, Open_32, 
            Open_33, Open_34, Open_35, Open_36, Open_37}), .ROM_DAT_O({ROM_DAT_O}), 
            .w_clk_cpu(w_clk_cpu), .n87({n87}), .\counter[2] (\counter[2] ), 
            .\LM32D_DAT_O[15] (LM32D_DAT_O[15]), .\SHAREDBUS_SEL_I[1] (\SHAREDBUS_SEL_I[1] ), 
            .n41490(n41490), .ROM_ACK_O(ROM_ACK_O), .n42726(n42726), .\data[21] (\data[21] ), 
            .\LM32D_DAT_O[14] (LM32D_DAT_O[14]), .\LM32D_DAT_O[13] (LM32D_DAT_O[13]), 
            .\LM32D_DAT_O[12] (LM32D_DAT_O[12]), .\LM32D_DAT_O[11] (LM32D_DAT_O[11]), 
            .\data[19] (\data[19] ), .\LM32D_DAT_O[10] (LM32D_DAT_O[10]), 
            .\LM32D_DAT_O[9] (LM32D_DAT_O[9]), .w_clk_cpu_enable_303(w_clk_cpu_enable_303), 
            .\data[30] (\data[30] ), .\LM32D_DAT_O[8] (LM32D_DAT_O[8]), 
            .\LM32D_DAT_O[7] (LM32D_DAT_O[7]), .n41426(n41426), .\LM32D_DAT_O[0] (LM32D_DAT_O[0]), 
            .\LM32D_DAT_O[6] (LM32D_DAT_O[6]), .\data[29] (\data[29] ), 
            .\data[28] (\data[28] ), .n93({n93}), .n92({n92}), .n41422(n41422), 
            .n41435(n41435), .n35(n35), .\data[27] (\data[27] ), .\data[26] (\data[26] ), 
            .\data[25] (\data[25] ), .\data[18] (\data[18] ), .\data[24] (\data[24] ), 
            .\LM32D_DAT_O[5] (LM32D_DAT_O[5]), .\LM32D_DAT_O[4] (LM32D_DAT_O[4]), 
            .\LM32D_DAT_O[3] (LM32D_DAT_O[3]), .\LM32D_DAT_O[2] (LM32D_DAT_O[2]), 
            .\data[23] (\data[23] ), .\LM32D_DAT_O[1] (LM32D_DAT_O[1]), 
            .\data[17] (\data[17] ), .\data[16] (\data[16] ), .n96({n96}), 
            .\data[22] (\data[22] ), .\data[20] (\data[20] ), .GND_net(GND_net), 
            .\SHAREDBUS_ADR_I[10] (\SHAREDBUS_ADR_I[10] ), .\SHAREDBUS_ADR_I[9] (\SHAREDBUS_ADR_I[9] ), 
            .\SHAREDBUS_ADR_I[8] (\SHAREDBUS_ADR_I[8] ), .\SHAREDBUS_ADR_I[7] (\SHAREDBUS_ADR_I[7] ), 
            .\SHAREDBUS_ADR_I[6] (\SHAREDBUS_ADR_I[6] ), .\SHAREDBUS_ADR_I[5] (\SHAREDBUS_ADR_I[5] ), 
            .\SHAREDBUS_ADR_I[4] (\SHAREDBUS_ADR_I[4] ), .\SHAREDBUS_ADR_I[3] (\SHAREDBUS_ADR_I[3] ), 
            .\SHAREDBUS_ADR_I[2] (\SHAREDBUS_ADR_I[2] ), .VCC_net(VCC_net), 
            .counter_2__N_178(counter_2__N_178)) /* synthesis syn_module_defined=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_top.v(398[17] 413[8])
    
endmodule
//
// Verilog Description of module jtag_cores
// module not written out since it is a black-box. 
//

//
// Verilog Description of module lm32_cpu
//

module lm32_cpu (w_result, w_clk_cpu, data_bus_error_exception_N_1225, 
            n42726, read_idx_0_d, n23059, n23091, n23058, n23090, 
            n23067, n23099, LM32D_CYC_O, n23068, n23100, LM32I_CYC_O, 
            n42734, n42738, read_idx_1_d, n23069, n23101, n42732, 
            n23070, n23102, n23071, n23103, n23072, n23104, \counter[2] , 
            n41470, write_idx_w, n23185, n23186, n23073, n23105, 
            n23074, n23106, n23075, n23107, n23076, n23108, n22885, 
            \jtag_reg_addr_d[0] , \jtag_reg_addr_d[1] , wb_load_complete_N_2129, 
            GND_net, reg_data_1, n23056, n23088, n23057, n23089, 
            n22999, n22877, n22874, n23053, n23085, n23054, n23086, 
            n23060, n23092, n23061, n23093, n23062, n23094, n23063, 
            n23095, n23064, n23096, n23065, n23097, n23066, n23098, 
            n23052, n23084, n23055, n23087, n23077, n23109, n23078, 
            n23110, n23079, n23111, n23080, n23112, n23081, n23113, 
            n23082, n23114, n23083, n23115, i_cyc_o_N_1759, LM32D_WE_O, 
            LM32D_DAT_O, SHAREDBUS_DAT_O, LM32D_ADR_O, LM32D_SEL_O, 
            LM32D_STB_O, jtag_reg_d, jtag_reg_q, jtag_update_N_2932, 
            jtag_reg_addr_q, \LM32I_ADR_O[2] , \selected_1__N_344[0] , 
            \LM32I_ADR_O[31] , bus_error_f_N_1764, \LM32I_ADR_O[30] , 
            \LM32I_ADR_O[29] , \LM32I_ADR_O[28] , \LM32I_ADR_O[27] , \LM32I_ADR_O[26] , 
            \LM32I_ADR_O[25] , \LM32I_ADR_O[24] , \LM32I_ADR_O[23] , \LM32I_ADR_O[22] , 
            \LM32I_ADR_O[21] , \LM32I_ADR_O[20] , \LM32I_ADR_O[19] , \LM32I_ADR_O[18] , 
            \LM32I_ADR_O[17] , \LM32I_ADR_O[16] , \LM32I_ADR_O[15] , \LM32I_ADR_O[14] , 
            \LM32I_ADR_O[13] , \LM32I_ADR_O[12] , \LM32I_ADR_O[11] , \LM32I_ADR_O[10] , 
            \LM32I_ADR_O[9] , \LM32I_ADR_O[8] , \LM32I_ADR_O[7] , \LM32I_ADR_O[6] , 
            \LM32I_ADR_O[5] , \LM32I_ADR_O[4] , \LM32I_ADR_O[3] , n41479, 
            n38871) /* synthesis syn_module_defined=1 */ ;
    output [31:0]w_result;
    input w_clk_cpu;
    input data_bus_error_exception_N_1225;
    input n42726;
    output [4:0]read_idx_0_d;
    input n23059;
    input n23091;
    input n23058;
    input n23090;
    input n23067;
    input n23099;
    output LM32D_CYC_O;
    input n23068;
    input n23100;
    output LM32I_CYC_O;
    output n42734;
    output n42738;
    output [4:0]read_idx_1_d;
    input n23069;
    input n23101;
    output n42732;
    input n23070;
    input n23102;
    input n23071;
    input n23103;
    input n23072;
    input n23104;
    input \counter[2] ;
    output n41470;
    output [4:0]write_idx_w;
    output n23185;
    output n23186;
    input n23073;
    input n23105;
    input n23074;
    input n23106;
    input n23075;
    input n23107;
    input n23076;
    input n23108;
    input n22885;
    output \jtag_reg_addr_d[0] ;
    output \jtag_reg_addr_d[1] ;
    input wb_load_complete_N_2129;
    input GND_net;
    input [31:0]reg_data_1;
    input n23056;
    input n23088;
    input n23057;
    input n23089;
    input n22999;
    output n22877;
    output n22874;
    input n23053;
    input n23085;
    input n23054;
    input n23086;
    input n23060;
    input n23092;
    input n23061;
    input n23093;
    input n23062;
    input n23094;
    input n23063;
    input n23095;
    input n23064;
    input n23096;
    input n23065;
    input n23097;
    input n23066;
    input n23098;
    input n23052;
    input n23084;
    input n23055;
    input n23087;
    input n23077;
    input n23109;
    input n23078;
    input n23110;
    input n23079;
    input n23111;
    input n23080;
    input n23112;
    input n23081;
    input n23113;
    input n23082;
    input n23114;
    input n23083;
    input n23115;
    input i_cyc_o_N_1759;
    output LM32D_WE_O;
    output [31:0]LM32D_DAT_O;
    input [31:0]SHAREDBUS_DAT_O;
    output [31:0]LM32D_ADR_O;
    output [3:0]LM32D_SEL_O;
    output LM32D_STB_O;
    output [7:0]jtag_reg_d;
    input [7:0]jtag_reg_q;
    input jtag_update_N_2932;
    input [2:0]jtag_reg_addr_q;
    output \LM32I_ADR_O[2] ;
    output \selected_1__N_344[0] ;
    output \LM32I_ADR_O[31] ;
    input bus_error_f_N_1764;
    output \LM32I_ADR_O[30] ;
    output \LM32I_ADR_O[29] ;
    output \LM32I_ADR_O[28] ;
    output \LM32I_ADR_O[27] ;
    output \LM32I_ADR_O[26] ;
    output \LM32I_ADR_O[25] ;
    output \LM32I_ADR_O[24] ;
    output \LM32I_ADR_O[23] ;
    output \LM32I_ADR_O[22] ;
    output \LM32I_ADR_O[21] ;
    output \LM32I_ADR_O[20] ;
    output \LM32I_ADR_O[19] ;
    output \LM32I_ADR_O[18] ;
    output \LM32I_ADR_O[17] ;
    output \LM32I_ADR_O[16] ;
    output \LM32I_ADR_O[15] ;
    output \LM32I_ADR_O[14] ;
    output \LM32I_ADR_O[13] ;
    output \LM32I_ADR_O[12] ;
    output \LM32I_ADR_O[11] ;
    output \LM32I_ADR_O[10] ;
    output \LM32I_ADR_O[9] ;
    output \LM32I_ADR_O[8] ;
    output \LM32I_ADR_O[7] ;
    output \LM32I_ADR_O[6] ;
    output \LM32I_ADR_O[5] ;
    output \LM32I_ADR_O[4] ;
    output \LM32I_ADR_O[3] ;
    input n41479;
    input n38871;
    
    wire w_clk_cpu /* synthesis SET_AS_NETWORK=w_clk_cpu, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(22[6:15])
    wire jtag_update_N_2932 /* synthesis is_inv_clock=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(203[14:23])
    wire [31:0]w_result_31__N_680;
    wire [31:0]load_data_w;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(679[23:34])
    
    wire w_result_sel_load_w, data_bus_error_exception, exception_m;
    wire [31:0]logic_result_x;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(566[23:37])
    wire [31:0]mc_result_x;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(616[23:34])
    
    wire x_result_sel_mc_arith_x;
    wire [31:0]n1253;
    wire [31:0]sext_result_x;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(572[23:36])
    
    wire x_result_sel_sext_x;
    wire [31:0]x_result_31__N_1066;
    
    wire n3, n7;
    wire [4:0]csr_x;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(478[22:27])
    
    wire n10;
    wire [31:2]branch_target_m;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(411[20:35])
    
    wire w_clk_cpu_enable_985, n22503;
    wire [31:2]branch_target_x;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(410[20:35])
    
    wire branch_taken_m, stall_a_N_1256, n4, n41199, n37259, w_clk_cpu_enable_984;
    wire [29:0]branch_target_x_31__N_1122;
    wire [31:0]n23116;
    wire [31:0]m_result;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(520[22:30])
    wire [31:0]operand_w_31__N_1187;
    
    wire n42746;
    wire [31:0]operand_w_31__N_840;
    wire [31:2]pc_m;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(634[21:25])
    wire [31:2]memop_pc_w;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(514[20:30])
    
    wire data_bus_error_exception_m, stall_a_N_1259, n41513, n41512;
    wire [31:0]operand_1_x;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(524[22:33])
    wire [31:0]d_result_1;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(518[22:32])
    
    wire n41526;
    wire [31:8]deba;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(732[28:32])
    
    wire n41540, n41428, branch_flushX_m_N_1116, n41408, csr_write_enable_x, 
        valid_x, n41365, valid_w, valid_m, n22501, n41466, x_result_sel_sext_N_1782, 
        x_result_sel_add_x, x_result_sel_add_N_1785, w_result_sel_load_m, 
        w_clk_cpu_enable_972, load_x, n3_adj_3776, n7_adj_3777, n10_adj_3778, 
        jtag_break, break_x, non_debug_exception_x_N_1357, n41430, m_bypass_enable_m, 
        x_bypass_enable_x, interlock_N_1333, interlock_N_1327, bus_error_x;
    wire [2:0]eid_x_2__N_1098;
    
    wire n31712, cycles_5__N_2495, n41395, n7_adj_3779, bret_x, bret_q_x, 
        n7_adj_3780, n7_adj_3781, n7_adj_3782, n7_adj_3783, n7_adj_3784, 
        n7_adj_3785, n7_adj_3786, n7_adj_3787, n7_adj_3788, n7_adj_3789, 
        n31636, n7_adj_3790, n7_adj_3791, n7_adj_3792, n7_adj_3793, 
        n7_adj_3794, n41391, n7_adj_3795, stall_wb_load, n52, n7_adj_3796, 
        n41576, n41577;
    wire [29:0]branch_target_m_31__N_1157;
    
    wire exception_m_N_1355, w_clk_cpu_enable_711, w_clk_cpu_enable_878, 
        n39086, n41573, n41574, n23901, n41530;
    wire [31:8]eba;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(730[28:31])
    
    wire n3_adj_3797, n3_adj_3798, n3_adj_3799, n3_adj_3800, n41444, 
        n41320, n41319, n41321, n3_adj_3801, n10_adj_3802, n3_adj_3803, 
        n3_adj_3804, n3_adj_3805, n3_adj_3806, n3_adj_3807, n3_adj_3808, 
        n3_adj_3809, n3_adj_3810;
    wire [31:2]branch_target_d;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(397[21:36])
    wire [31:0]bypass_data_0;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(543[22:35])
    
    wire n22224, n3_adj_3811, n3_adj_3812, n3_adj_3813, n3_adj_3814, 
        n3_adj_3815, n3_adj_3816, write_enable_w, n41531, dc_re, n41544, 
        n41570, n41571, n41543, n36634;
    wire [31:2]pc_d;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(632[21:25])
    wire [31:0]instruction_d;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(654[30:43])
    
    wire valid_f, valid_f_N_1227, n39126;
    wire [31:0]store_operand_x;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(525[22:37])
    wire [31:0]bypass_data_1;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(544[22:35])
    
    wire eba_31__N_1101;
    wire [31:0]muliplicand;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(90[22:33])
    
    wire n36633, n41547;
    wire [31:0]operand_w;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(527[22:31])
    wire [4:0]write_idx_m;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(475[25:36])
    
    wire w_result_sel_mul_w, w_result_sel_mul_m, deba_31__N_1120, write_enable_m, 
        debug_exception_w, debug_exception_m, non_debug_exception_w, non_debug_exception_m, 
        n10_adj_3817, n36632, n41567, n41568;
    wire [31:0]adder_result_x;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(559[23:37])
    wire [31:0]x_result_31__N_616;
    
    wire n10_adj_3818, m_result_sel_compare_x, n41419, n10_adj_3819, 
        n41147, n38972, n25563, n41564, n41565, n36631;
    wire [4:0]write_idx_x;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(474[25:36])
    
    wire n26142;
    wire [4:0]write_idx_4__N_1770;
    
    wire m_result_sel_shift_m, m_result_sel_shift_x, n41561, n41562, 
        memop_pc_w_31__N_1219, m_result_sel_compare_m, n24298, n1, n2, 
        n41361, w_clk_cpu_enable_697, n1_adj_3820, n2_adj_3821, n29325;
    wire [31:0]im;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(141[22:24])
    
    wire n36690, n38878;
    wire [31:0]csr_read_data_x;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(628[22:37])
    
    wire n1_adj_3822, n2_adj_3823, x_result_sel_csr_x, branch_m, n39497;
    wire [31:0]x_result;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(519[22:30])
    
    wire raw_x_0;
    wire [31:0]bypass_data_0_31__N_872;
    
    wire raw_w_0;
    wire [31:0]bypass_data_0_31__N_1002;
    
    wire n1_adj_3824, n2_adj_3825, n1_adj_3826, n2_adj_3827, n1_adj_3828, 
        n2_adj_3829, n1_adj_3830, n2_adj_3831, n27, n1_adj_3832, n2_adj_3833, 
        n26, n22, n10_adj_3834, n20, n41546, n1_adj_3835, n2_adj_3836, 
        n41451, n41372, n26096, n1_adj_3837, n2_adj_3838, w_clk_cpu_enable_245, 
        n1_adj_3839, n2_adj_3840;
    wire [31:0]n21231;
    
    wire n9, n39068, n41503, n1_adj_3841, n2_adj_3842, n36630, n38764, 
        n41411, n1_adj_3843, n2_adj_3844;
    wire [31:0]jrx_csr_read_data;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(686[23:40])
    
    wire raw_x_1, n39329, n10_adj_3845, n4_adj_3846, n1_adj_3847, 
        n2_adj_3848, n10_adj_3849, n31, n1_adj_3850, n2_adj_3851, 
        n1_adj_3852, n2_adj_3853, n10_adj_3854, n36629, n41375, n39970, 
        n1_adj_3855, n2_adj_3856, n1_adj_3857, n2_adj_3858, n10_adj_3859, 
        n10_adj_3860, scall_x, scall_d, n1_adj_3861, n2_adj_3862, 
        n1_adj_3863, n2_adj_3864, n1_adj_3865, n2_adj_3866, n1_adj_3867, 
        n2_adj_3868, n1_adj_3869, n2_adj_3870, n41555, n41556, n10_adj_3871, 
        n36628, n1_adj_3872, n2_adj_3873, n40567, n1_adj_3874, n2_adj_3875, 
        n1_adj_3876, n2_adj_3877, n1_adj_3878, n2_adj_3879, n1_adj_3880, 
        n36772;
    wire [31:0]multiplier_result_w;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(597[23:42])
    
    wire n10_adj_3881, n1_adj_3882, n2_adj_3883, condition_met_m, n41507, 
        n1_adj_3884, n2_adj_3885, n1_adj_3886, n2_adj_3887, n1_adj_3888, 
        n2_adj_3889, n10_adj_3890, n10_adj_3891, n41552, n41553, n36493, 
        cmp_zero, n36627, n9_adj_3892, n7_adj_3893, n8;
    wire [31:0]bypass_data_1_31__N_1034;
    wire [31:0]bypass_data_1_31__N_904;
    
    wire n36626, n10_adj_3894, n41549, n41550, n10_adj_3895, n10_adj_3896;
    wire [31:0]operand_m;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(526[22:31])
    wire [31:0]m_result_31__N_648;
    
    wire n40566, n40565, n10_adj_3897, n39056, n23668, n39064, n18863, 
        branch_x, branch_d;
    wire [4:0]write_idx_m_4__N_1152;
    
    wire valid_d, n41387, n25722, n41373;
    wire [4:0]write_idx_d;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(473[26:37])
    
    wire write_enable_x, n25724, n38799;
    wire [2:0]condition_x;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(480[27:38])
    wire [1:0]size_x;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(392[22:28])
    
    wire n41491;
    wire [3:0]byte_enable_x;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(245[29:42])
    
    wire n41492, n41580, n41579, load_m, wb_select_m, wb_load_complete, 
        n41493, n41583, n39775, n39776;
    wire [3:0]logic_op_x;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(565[26:36])
    
    wire condition_met_x, n41582, n41586, n41585;
    wire [3:0]logic_op_d;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(564[27:37])
    
    wire n39363, n41589;
    wire [31:0]instruction;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(195[31:42])
    
    wire n41588;
    wire [1:0]size_d;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(391[23:29])
    
    wire n41592, n46, w_clk_cpu_enable_886, n41591, n36625, n41595, 
        n41594, n41598, n41597, n41601, raw_w_1, n41600, n41604, 
        n41603, n41607, n41606, n41610, n41609, n25705, n41359, 
        n41613, n18869, n41612;
    wire [2:0]eid_x_2__N_999;
    
    wire reset_exception, store_x, n42730, n42736;
    wire [31:0]shifter_result_m;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(583[23:39])
    
    wire n23893, n38801, n36624, n36623, n39459, n34433, n39886, 
        n6, n39890, n36488, n36489, n36492, n36487, n36622, n36621, 
        n41438;
    wire [31:0]left_shift_result;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(93[22:39])
    wire [31:0]n1826;
    
    wire n42722, n41397, n39334, n36491, branch_predict_m, branch_predict_taken_m, 
        eret_x, n4_adj_3898, eie, ie_N_2822, ie_N_2821, jtag_reg_d_7__N_505, 
        w_clk_cpu_enable_638, valid_d_N_1264, n36490, n22524, write_enable_m_N_1313, 
        w_clk_cpu_enable_958, n38840, n41502, n41394, n41457, n41504, 
        n36486, m_result_sel_shift_d, w_result_sel_mul_x, w_result_sel_mul_d, 
        x_bypass_enable_d, n41459, m_bypass_enable_x, m_bypass_enable_d;
    wire [23:0]n21411;
    
    wire adder_carry_n_x, write_enable_N_1809, adder_op_x_n, adder_op_d_N_1339, 
        branch_predict_x, branch_predict_d, branch_predict_taken_x, mc_stall_request_x, 
        divide_by_zero_x, n31661, n26126, eret_d, bret_d, bus_error_d, 
        n41406, n40464, store_d, n41432, adder_op_x, n41376, n41541, 
        store_m, n4_adj_3899, n41474, n9_adj_3900, n24748, n39150, 
        n3_adj_3901, n39082, n38827, n4_adj_3902, raw_m_0, n41472, 
        ie, bie_N_2835, n25625, n41351, n39892, n39222, n2_adj_3903, 
        n41473, n23750, n39142, n2_adj_3904;
    wire [31:0]store_data_x;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(243[22:34])
    
    wire n36706, n2_adj_3905, n36708, bie, dc_re_N_2934, n30, n29, 
        break_d, direction_x, sign_extend_x, n41384, x_result_sel_csr_d, 
        direction_m, w_clk_cpu_enable_623, n26122;
    wire [31:0]d_result_0;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(517[22:32])
    
    wire n18875, n41417, w_clk_cpu_enable_865, n41364, n22236, n41380, 
        sign_extend_immediate, n41367, n13, n41407;
    wire [31:2]pc_f;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(631[21:25])
    
    wire n42740, w_clk_cpu_enable_216, n37179, n41345;
    wire [31:0]n1760;
    
    wire stall_wb_load_N_2112, w_clk_cpu_enable_914, n41357, w_clk_cpu_enable_763, 
        w_clk_cpu_enable_330, w_clk_cpu_enable_983, n38725;
    
    PFUMX w_result_31__I_0_i3 (.BLUT(w_result_31__N_680[2]), .ALUT(load_data_w[2]), 
          .C0(w_result_sel_load_w), .Z(w_result[2])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3IX data_bus_error_seen_616 (.D(n42726), .SP(data_bus_error_exception_N_1225), 
            .CD(exception_m), .CK(w_clk_cpu), .Q(data_bus_error_exception));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2200[5] 2207[8])
    defparam data_bus_error_seen_616.GSR = "ENABLED";
    PFUMX w_result_31__I_0_i4 (.BLUT(w_result_31__N_680[3]), .ALUT(load_data_w[3]), 
          .C0(w_result_sel_load_w), .Z(w_result[3])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i5 (.BLUT(w_result_31__N_680[4]), .ALUT(load_data_w[4]), 
          .C0(w_result_sel_load_w), .Z(w_result[4])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_75_i28_3_lut (.A(logic_result_x[27]), .B(mc_result_x[27]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i28_3_lut.init = 16'hcaca;
    LUT4 mux_76_i32_3_lut (.A(n1253[31]), .B(sext_result_x[15]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i32_3_lut.init = 16'hcaca;
    LUT4 mux_76_i31_3_lut (.A(n1253[30]), .B(sext_result_x[15]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i31_3_lut.init = 16'hcaca;
    PFUMX i23 (.BLUT(n3), .ALUT(n7), .C0(csr_x[3]), .Z(n10));
    FD1P3IX branch_target_m_i2_i3 (.D(branch_target_x[3]), .SP(w_clk_cpu_enable_985), 
            .CD(n22503), .CK(w_clk_cpu), .Q(branch_target_m[3])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i3.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(branch_taken_m), .B(stall_a_N_1256), .C(n4), .D(n41199), 
         .Z(n37259)) /* synthesis lut_function=(!(A+!(B (C+(D))+!B (C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1890[6] 1900[7])
    defparam i1_4_lut.init = 16'h5450;
    PFUMX w_result_31__I_0_i6 (.BLUT(w_result_31__N_680[5]), .ALUT(load_data_w[5]), 
          .C0(w_result_sel_load_w), .Z(w_result[5])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_76_i30_3_lut (.A(n1253[29]), .B(sext_result_x[15]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i30_3_lut.init = 16'hcaca;
    LUT4 mux_76_i29_3_lut (.A(n1253[28]), .B(sext_result_x[15]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i29_3_lut.init = 16'hcaca;
    FD1P3AX csr_x_i0_i1 (.D(read_idx_0_d[1]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(csr_x[1])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam csr_x_i0_i1.GSR = "ENABLED";
    FD1P3AX branch_target_x_i2_i31 (.D(branch_target_x_31__N_1122[29]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[31])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i31.GSR = "ENABLED";
    LUT4 mux_76_i28_3_lut (.A(n1253[27]), .B(sext_result_x[15]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i28_3_lut.init = 16'hcaca;
    LUT4 mux_20532_i8_3_lut (.A(n23059), .B(n23091), .C(read_idx_0_d[4]), 
         .Z(n23116[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i8_3_lut.init = 16'hcaca;
    LUT4 mux_20532_i7_3_lut (.A(n23058), .B(n23090), .C(read_idx_0_d[4]), 
         .Z(n23116[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i7_3_lut.init = 16'hcaca;
    LUT4 mux_20532_i16_3_lut (.A(n23067), .B(n23099), .C(read_idx_0_d[4]), 
         .Z(n23116[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i16_3_lut.init = 16'hcaca;
    LUT4 m_result_31__I_0_i16_3_lut (.A(m_result[15]), .B(operand_w_31__N_1187[15]), 
         .C(n42746), .Z(operand_w_31__N_840[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i16_3_lut.init = 16'hcaca;
    LUT4 mux_19174_i14_3_lut (.A(pc_m[15]), .B(memop_pc_w[15]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i14_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut (.A(LM32D_CYC_O), .B(stall_a_N_1259), .C(n41513), .D(n41512), 
         .Z(stall_a_N_1256)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(746[5:16])
    defparam i2_4_lut.init = 16'hfeee;
    FD1P3AX operand_1_x_i0_i14 (.D(d_result_1[14]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[14])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i14.GSR = "ENABLED";
    FD1P3AX operand_1_x_i0_i13 (.D(d_result_1[13]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[13])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i13.GSR = "ENABLED";
    FD1P3AX operand_1_x_i0_i12 (.D(d_result_1[12]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[12])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i12.GSR = "ENABLED";
    FD1P3AX operand_1_x_i0_i11 (.D(d_result_1[11]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[11])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i11.GSR = "ENABLED";
    FD1P3AX operand_1_x_i0_i10 (.D(d_result_1[10]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[10])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i10.GSR = "ENABLED";
    LUT4 mux_76_i27_3_lut (.A(n1253[26]), .B(sext_result_x[15]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i27_3_lut.init = 16'hcaca;
    FD1P3AX operand_1_x_i0_i9 (.D(d_result_1[9]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[9])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i9.GSR = "ENABLED";
    FD1P3AX operand_1_x_i0_i8 (.D(d_result_1[8]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[8])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i8.GSR = "ENABLED";
    FD1P3AX operand_1_x_i0_i7 (.D(d_result_1[7]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[7])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i7.GSR = "ENABLED";
    FD1P3AX operand_1_x_i0_i6 (.D(d_result_1[6]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[6])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i6.GSR = "ENABLED";
    FD1P3AX operand_1_x_i0_i5 (.D(d_result_1[5]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[5])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i5.GSR = "ENABLED";
    FD1P3AX operand_1_x_i0_i4 (.D(d_result_1[4]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[4])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i4.GSR = "ENABLED";
    FD1P3AX operand_1_x_i0_i3 (.D(d_result_1[3]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[3])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i3.GSR = "ENABLED";
    LUT4 mux_465_i7_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[8]), .C(branch_target_x[8]), 
         .Z(n41540)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i7_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    FD1P3AX operand_1_x_i0_i2 (.D(d_result_1[2]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[2])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i2.GSR = "ENABLED";
    FD1P3AX operand_1_x_i0_i1 (.D(d_result_1[1]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[1])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i1.GSR = "ENABLED";
    LUT4 branch_flushX_m_I_0_700_2_lut_rep_321 (.A(n41428), .B(branch_flushX_m_N_1116), 
         .Z(n41408)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1676[29] 1687[9])
    defparam branch_flushX_m_I_0_700_2_lut_rep_321.init = 16'h4444;
    LUT4 mux_76_i26_3_lut (.A(n1253[25]), .B(sext_result_x[15]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i26_3_lut.init = 16'hcaca;
    FD1P3AX branch_target_x_i2_i30 (.D(branch_target_x_31__N_1122[28]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[30])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i30.GSR = "ENABLED";
    FD1P3AX branch_target_x_i2_i29 (.D(branch_target_x_31__N_1122[27]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[29])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i29.GSR = "ENABLED";
    PFUMX w_result_31__I_0_i7 (.BLUT(w_result_31__N_680[6]), .ALUT(load_data_w[6]), 
          .C0(w_result_sel_load_w), .Z(w_result[6])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 csr_write_enable_x_I_0_2_lut_rep_278_3_lut_4_lut (.A(n41428), .B(branch_flushX_m_N_1116), 
         .C(csr_write_enable_x), .D(valid_x), .Z(n41365)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1676[29] 1687[9])
    defparam csr_write_enable_x_I_0_2_lut_rep_278_3_lut_4_lut.init = 16'hb000;
    LUT4 m_result_31__I_0_i15_3_lut (.A(m_result[14]), .B(operand_w_31__N_1187[14]), 
         .C(n42746), .Z(operand_w_31__N_840[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i15_3_lut.init = 16'hcaca;
    LUT4 mux_19174_i13_3_lut (.A(pc_m[14]), .B(memop_pc_w[14]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i13_3_lut.init = 16'hcaca;
    FD1P3AX branch_target_x_i2_i28 (.D(branch_target_x_31__N_1122[26]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[28])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i28.GSR = "ENABLED";
    FD1P3AX branch_target_x_i2_i27 (.D(branch_target_x_31__N_1122[25]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[27])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i27.GSR = "ENABLED";
    FD1S3IX valid_w_621 (.D(valid_m), .CK(w_clk_cpu), .CD(n41428), .Q(valid_w));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2264[5] 2299[8])
    defparam valid_w_621.GSR = "ENABLED";
    FD1P3IX x_result_sel_mc_arith_x_627 (.D(n41466), .SP(w_clk_cpu_enable_984), 
            .CD(n22501), .CK(w_clk_cpu), .Q(x_result_sel_mc_arith_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam x_result_sel_mc_arith_x_627.GSR = "ENABLED";
    FD1P3IX x_result_sel_sext_x_628 (.D(x_result_sel_sext_N_1782), .SP(w_clk_cpu_enable_984), 
            .CD(n22501), .CK(w_clk_cpu), .Q(x_result_sel_sext_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam x_result_sel_sext_x_628.GSR = "ENABLED";
    FD1P3IX x_result_sel_add_x_630 (.D(x_result_sel_add_N_1785), .SP(w_clk_cpu_enable_984), 
            .CD(n22501), .CK(w_clk_cpu), .Q(x_result_sel_add_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam x_result_sel_add_x_630.GSR = "ENABLED";
    FD1P3IX w_result_sel_load_m_663 (.D(load_x), .SP(w_clk_cpu_enable_972), 
            .CD(n22503), .CK(w_clk_cpu), .Q(w_result_sel_load_m));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam w_result_sel_load_m_663.GSR = "ENABLED";
    FD1P3AX branch_target_x_i2_i26 (.D(branch_target_x_31__N_1122[24]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[26])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i26.GSR = "ENABLED";
    FD1P3AX branch_target_x_i2_i25 (.D(branch_target_x_31__N_1122[23]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[25])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i25.GSR = "ENABLED";
    PFUMX i23_adj_275 (.BLUT(n3_adj_3776), .ALUT(n7_adj_3777), .C0(csr_x[3]), 
          .Z(n10_adj_3778));
    LUT4 breakpoint_exception_I_56_3_lut_rep_439 (.A(valid_x), .B(jtag_break), 
         .C(break_x), .Z(n41526)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam breakpoint_exception_I_56_3_lut_rep_439.init = 16'hecec;
    LUT4 i1_2_lut_rep_343_4_lut (.A(valid_x), .B(jtag_break), .C(break_x), 
         .D(non_debug_exception_x_N_1357), .Z(n41430)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam i1_2_lut_rep_343_4_lut.init = 16'hffec;
    LUT4 i1_4_lut_adj_276 (.A(m_bypass_enable_m), .B(x_bypass_enable_x), 
         .C(interlock_N_1333), .D(interlock_N_1327), .Z(n4)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (C+(D))))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1890[6] 1900[7])
    defparam i1_4_lut_adj_276.init = 16'h7350;
    FD1P3AX operand_1_x_i0_i0 (.D(d_result_1[0]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[0])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i0.GSR = "ENABLED";
    LUT4 mux_76_i25_3_lut (.A(n1253[24]), .B(sext_result_x[15]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i25_3_lut.init = 16'hcaca;
    LUT4 i28947_2_lut_3_lut_4_lut (.A(valid_x), .B(jtag_break), .C(break_x), 
         .D(bus_error_x), .Z(eid_x_2__N_1098[0])) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam i28947_2_lut_3_lut_4_lut.init = 16'hfdff;
    LUT4 m_result_31__I_0_i14_3_lut (.A(m_result[13]), .B(operand_w_31__N_1187[13]), 
         .C(n42746), .Z(operand_w_31__N_840[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i14_3_lut.init = 16'hcaca;
    LUT4 i29151_2_lut_2_lut_3_lut_4_lut (.A(csr_x[2]), .B(csr_x[1]), .C(csr_x[4]), 
         .D(csr_x[3]), .Z(n31712)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i29151_2_lut_2_lut_3_lut_4_lut.init = 16'hfeff;
    LUT4 i28948_2_lut_rep_308_3_lut (.A(n41428), .B(branch_flushX_m_N_1116), 
         .C(cycles_5__N_2495), .Z(n41395)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1676[29] 1687[9])
    defparam i28948_2_lut_rep_308_3_lut.init = 16'hf4f4;
    FD1P3AX branch_target_x_i2_i24 (.D(branch_target_x_31__N_1122[22]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[24])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i24.GSR = "ENABLED";
    FD1P3AX branch_target_x_i2_i23 (.D(branch_target_x_31__N_1122[21]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[23])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i23.GSR = "ENABLED";
    LUT4 i2_2_lut_3_lut (.A(csr_x[2]), .B(csr_x[1]), .C(deba[9]), .Z(n7_adj_3779)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut.init = 16'h1010;
    LUT4 i2_2_lut_3_lut_adj_277 (.A(csr_x[2]), .B(csr_x[1]), .C(deba[26]), 
         .Z(n7_adj_3777)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut_adj_277.init = 16'h1010;
    LUT4 mux_19174_i12_3_lut (.A(pc_m[13]), .B(memop_pc_w[13]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i12_3_lut.init = 16'hcaca;
    LUT4 mux_20532_i17_3_lut (.A(n23068), .B(n23100), .C(read_idx_0_d[4]), 
         .Z(n23116[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i17_3_lut.init = 16'hcaca;
    PFUMX w_result_31__I_0_i8 (.BLUT(w_result_31__N_680[7]), .ALUT(load_data_w[7]), 
          .C0(w_result_sel_load_w), .Z(w_result[7])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 bret_x_I_0_2_lut_3_lut_4_lut (.A(n41428), .B(branch_flushX_m_N_1116), 
         .C(bret_x), .D(valid_x), .Z(bret_q_x)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1676[29] 1687[9])
    defparam bret_x_I_0_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 i2_2_lut_3_lut_adj_278 (.A(csr_x[2]), .B(csr_x[1]), .C(deba[13]), 
         .Z(n7_adj_3780)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut_adj_278.init = 16'h1010;
    LUT4 i2_2_lut_3_lut_adj_279 (.A(csr_x[2]), .B(csr_x[1]), .C(deba[10]), 
         .Z(n7_adj_3781)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut_adj_279.init = 16'h1010;
    LUT4 i2_2_lut_3_lut_adj_280 (.A(csr_x[2]), .B(csr_x[1]), .C(deba[30]), 
         .Z(n7_adj_3782)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut_adj_280.init = 16'h1010;
    LUT4 mux_76_i24_3_lut (.A(n1253[23]), .B(sext_result_x[15]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i24_3_lut.init = 16'hcaca;
    FD1P3AX branch_target_x_i2_i22 (.D(branch_target_x_31__N_1122[20]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[22])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i22.GSR = "ENABLED";
    FD1P3AX branch_target_x_i2_i21 (.D(branch_target_x_31__N_1122[19]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[21])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i21.GSR = "ENABLED";
    LUT4 i2_2_lut_3_lut_adj_281 (.A(csr_x[2]), .B(csr_x[1]), .C(deba[12]), 
         .Z(n7_adj_3783)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut_adj_281.init = 16'h1010;
    LUT4 i2_2_lut_3_lut_adj_282 (.A(csr_x[2]), .B(csr_x[1]), .C(deba[16]), 
         .Z(n7_adj_3784)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut_adj_282.init = 16'h1010;
    LUT4 i2_2_lut_3_lut_adj_283 (.A(csr_x[2]), .B(csr_x[1]), .C(deba[23]), 
         .Z(n7_adj_3785)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut_adj_283.init = 16'h1010;
    LUT4 i2_2_lut_3_lut_adj_284 (.A(csr_x[2]), .B(csr_x[1]), .C(deba[19]), 
         .Z(n7_adj_3786)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut_adj_284.init = 16'h1010;
    LUT4 i2_2_lut_3_lut_adj_285 (.A(csr_x[2]), .B(csr_x[1]), .C(deba[15]), 
         .Z(n7_adj_3787)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut_adj_285.init = 16'h1010;
    LUT4 i2_2_lut_3_lut_adj_286 (.A(csr_x[2]), .B(csr_x[1]), .C(deba[22]), 
         .Z(n7_adj_3788)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut_adj_286.init = 16'h1010;
    LUT4 i2_2_lut_3_lut_adj_287 (.A(csr_x[2]), .B(csr_x[1]), .C(deba[21]), 
         .Z(n7_adj_3789)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut_adj_287.init = 16'h1010;
    PFUMX w_result_31__I_0_i9 (.BLUT(w_result_31__N_680[8]), .ALUT(load_data_w[8]), 
          .C0(w_result_sel_load_w), .Z(w_result[8])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i37929_2_lut_3_lut_3_lut_3_lut (.A(n41428), .B(branch_flushX_m_N_1116), 
         .C(cycles_5__N_2495), .Z(n31636)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1676[29] 1687[9])
    defparam i37929_2_lut_3_lut_3_lut_3_lut.init = 16'h0101;
    LUT4 i2_2_lut_3_lut_adj_288 (.A(csr_x[2]), .B(csr_x[1]), .C(deba[18]), 
         .Z(n7_adj_3790)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut_adj_288.init = 16'h1010;
    LUT4 m_result_31__I_0_i13_3_lut (.A(m_result[12]), .B(operand_w_31__N_1187[12]), 
         .C(n42746), .Z(operand_w_31__N_840[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i13_3_lut.init = 16'hcaca;
    LUT4 mux_19174_i11_3_lut (.A(pc_m[12]), .B(memop_pc_w[12]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i11_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_3_lut_adj_289 (.A(csr_x[2]), .B(csr_x[1]), .C(deba[14]), 
         .Z(n7_adj_3791)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut_adj_289.init = 16'h1010;
    LUT4 i2_2_lut_3_lut_adj_290 (.A(csr_x[2]), .B(csr_x[1]), .C(deba[25]), 
         .Z(n7_adj_3792)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut_adj_290.init = 16'h1010;
    FD1P3AX branch_target_x_i2_i20 (.D(branch_target_x_31__N_1122[18]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[20])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i20.GSR = "ENABLED";
    FD1P3AX branch_target_x_i2_i19 (.D(branch_target_x_31__N_1122[17]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[19])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i19.GSR = "ENABLED";
    LUT4 m_result_31__I_0_i12_3_lut (.A(m_result[11]), .B(operand_w_31__N_1187[11]), 
         .C(n42746), .Z(operand_w_31__N_840[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 mux_19174_i10_3_lut (.A(pc_m[11]), .B(memop_pc_w[11]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i10_3_lut.init = 16'hcaca;
    LUT4 mux_76_i23_3_lut (.A(n1253[22]), .B(sext_result_x[15]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i23_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_3_lut_adj_291 (.A(csr_x[2]), .B(csr_x[1]), .C(deba[28]), 
         .Z(n7_adj_3793)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut_adj_291.init = 16'h1010;
    LUT4 i2_2_lut_3_lut_adj_292 (.A(csr_x[2]), .B(csr_x[1]), .C(deba[24]), 
         .Z(n7_adj_3794)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut_adj_292.init = 16'h1010;
    LUT4 valid_x_I_0_2_lut_rep_304_3_lut (.A(n41428), .B(branch_flushX_m_N_1116), 
         .C(valid_x), .Z(n41391)) /* synthesis lut_function=(A (C)+!A !(B+!(C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1676[29] 1687[9])
    defparam valid_x_I_0_2_lut_rep_304_3_lut.init = 16'hb0b0;
    LUT4 i2_2_lut_3_lut_adj_293 (.A(csr_x[2]), .B(csr_x[1]), .C(deba[20]), 
         .Z(n7_adj_3795)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut_adj_293.init = 16'h1010;
    LUT4 i2_2_lut_3_lut_adj_294 (.A(csr_x[2]), .B(csr_x[1]), .C(deba[29]), 
         .Z(n7)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut_adj_294.init = 16'h1010;
    PFUMX w_result_31__I_0_i10 (.BLUT(w_result_31__N_680[9]), .ALUT(load_data_w[9]), 
          .C0(w_result_sel_load_w), .Z(w_result[9])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX branch_target_x_i2_i18 (.D(branch_target_x_31__N_1122[16]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[18])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i18.GSR = "ENABLED";
    FD1P3AX branch_target_x_i2_i17 (.D(branch_target_x_31__N_1122[15]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[17])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i17.GSR = "ENABLED";
    LUT4 stall_m_I_0_1_lut_rep_462 (.A(LM32I_CYC_O), .B(LM32D_CYC_O), .C(stall_wb_load), 
         .D(n52), .Z(w_clk_cpu_enable_972)) /* synthesis lut_function=(!(A+(B (C+(D))+!B (C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1924[21] 1957[39])
    defparam stall_m_I_0_1_lut_rep_462.init = 16'h0105;
    LUT4 mux_76_i22_3_lut (.A(n1253[21]), .B(sext_result_x[15]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i22_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_3_lut_adj_295 (.A(csr_x[2]), .B(csr_x[1]), .C(deba[31]), 
         .Z(n7_adj_3796)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut_adj_295.init = 16'h1010;
    PFUMX w_result_31__I_0_i11 (.BLUT(w_result_31__N_680[10]), .ALUT(load_data_w[10]), 
          .C0(w_result_sel_load_w), .Z(w_result[10])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_75_i29_3_lut (.A(logic_result_x[28]), .B(mc_result_x[28]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i29_3_lut.init = 16'hcaca;
    PFUMX i38595 (.BLUT(n41576), .ALUT(n41577), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[18]));
    LUT4 exception_x_I_0_2_lut_3_lut_4_lut (.A(n41428), .B(branch_flushX_m_N_1116), 
         .C(n41430), .D(valid_x), .Z(exception_m_N_1355)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1676[29] 1687[9])
    defparam exception_x_I_0_2_lut_3_lut_4_lut.init = 16'hb000;
    LUT4 stall_m_I_0_1_lut_rep_463 (.A(LM32I_CYC_O), .B(LM32D_CYC_O), .C(stall_wb_load), 
         .D(n52), .Z(w_clk_cpu_enable_711)) /* synthesis lut_function=(!(A+(B (C+(D))+!B (C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1924[21] 1957[39])
    defparam stall_m_I_0_1_lut_rep_463.init = 16'h0105;
    FD1P3AX branch_target_x_i2_i16 (.D(branch_target_x_31__N_1122[14]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[16])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i16.GSR = "ENABLED";
    FD1P3AX branch_target_x_i2_i15 (.D(branch_target_x_31__N_1122[13]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[15])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i15.GSR = "ENABLED";
    LUT4 mux_76_i21_3_lut (.A(n1253[20]), .B(sext_result_x[15]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i21_3_lut.init = 16'hcaca;
    LUT4 stall_m_I_0_1_lut_rep_464 (.A(LM32I_CYC_O), .B(LM32D_CYC_O), .C(stall_wb_load), 
         .D(n52), .Z(w_clk_cpu_enable_878)) /* synthesis lut_function=(!(A+(B (C+(D))+!B (C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1924[21] 1957[39])
    defparam stall_m_I_0_1_lut_rep_464.init = 16'h0105;
    LUT4 i36539_4_lut (.A(n42734), .B(n42738), .C(read_idx_1_d[3]), .D(read_idx_1_d[0]), 
         .Z(n39086)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i36539_4_lut.init = 16'h7bde;
    PFUMX i38593 (.BLUT(n41573), .ALUT(n41574), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[29]));
    LUT4 mux_76_i20_3_lut (.A(n1253[19]), .B(sext_result_x[15]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i20_3_lut.init = 16'hcaca;
    LUT4 i29120_2_lut_3_lut_3_lut_4_lut (.A(n41428), .B(branch_flushX_m_N_1116), 
         .C(valid_x), .D(cycles_5__N_2495), .Z(n23901)) /* synthesis lut_function=(A (C (D))+!A !(B+!(C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1676[29] 1687[9])
    defparam i29120_2_lut_3_lut_3_lut_4_lut.init = 16'hb000;
    FD1P3AX branch_target_x_i2_i14 (.D(branch_target_x_31__N_1122[12]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[14])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i14.GSR = "ENABLED";
    FD1P3AX branch_target_x_i2_i13 (.D(branch_target_x_31__N_1122[11]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[13])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i13.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_443 (.A(csr_x[2]), .B(csr_x[1]), .Z(n41530)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_443.init = 16'h8888;
    LUT4 i2_2_lut_3_lut_adj_296 (.A(csr_x[2]), .B(csr_x[1]), .C(eba[20]), 
         .Z(n3_adj_3797)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut_adj_296.init = 16'h8080;
    LUT4 i2_2_lut_3_lut_adj_297 (.A(csr_x[2]), .B(csr_x[1]), .C(eba[21]), 
         .Z(n3_adj_3798)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut_adj_297.init = 16'h8080;
    LUT4 i2_2_lut_3_lut_adj_298 (.A(csr_x[2]), .B(csr_x[1]), .C(eba[24]), 
         .Z(n3_adj_3799)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut_adj_298.init = 16'h8080;
    PFUMX w_result_31__I_0_i12 (.BLUT(w_result_31__N_680[11]), .ALUT(load_data_w[11]), 
          .C0(w_result_sel_load_w), .Z(w_result[11])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i2_2_lut_3_lut_adj_299 (.A(csr_x[2]), .B(csr_x[1]), .C(eba[28]), 
         .Z(n3_adj_3800)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut_adj_299.init = 16'h8080;
    LUT4 i2_3_lut_rep_357_4_lut (.A(csr_x[2]), .B(csr_x[1]), .C(csr_x[4]), 
         .D(csr_x[3]), .Z(n41444)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i2_3_lut_rep_357_4_lut.init = 16'h0800;
    LUT4 mux_20532_i18_3_lut (.A(n23069), .B(n23101), .C(read_idx_0_d[4]), 
         .Z(n23116[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i18_3_lut.init = 16'hcaca;
    PFUMX i38549 (.BLUT(n41320), .ALUT(n41319), .C0(csr_x[2]), .Z(n41321));
    PFUMX i23_adj_300 (.BLUT(n3_adj_3801), .ALUT(n7_adj_3788), .C0(csr_x[3]), 
          .Z(n10_adj_3802));
    LUT4 i2_2_lut_3_lut_adj_301 (.A(csr_x[2]), .B(csr_x[1]), .C(eba[22]), 
         .Z(n3_adj_3801)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut_adj_301.init = 16'h8080;
    LUT4 m_result_31__I_0_i11_3_lut (.A(m_result[10]), .B(operand_w_31__N_1187[10]), 
         .C(n42746), .Z(operand_w_31__N_840[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 mux_19174_i9_3_lut (.A(pc_m[10]), .B(memop_pc_w[10]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i9_3_lut.init = 16'hcaca;
    LUT4 m_result_31__I_0_i10_3_lut (.A(m_result[9]), .B(operand_w_31__N_1187[9]), 
         .C(n42746), .Z(operand_w_31__N_840[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i10_3_lut.init = 16'hcaca;
    LUT4 mux_19174_i8_3_lut (.A(pc_m[9]), .B(memop_pc_w[9]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i8_3_lut.init = 16'hcaca;
    LUT4 mux_76_i19_3_lut (.A(n1253[18]), .B(sext_result_x[15]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i19_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_3_lut_adj_302 (.A(csr_x[2]), .B(csr_x[1]), .C(eba[13]), 
         .Z(n3_adj_3803)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut_adj_302.init = 16'h8080;
    FD1P3AX branch_target_x_i2_i12 (.D(branch_target_x_31__N_1122[10]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[12])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i12.GSR = "ENABLED";
    FD1P3AX branch_target_x_i2_i11 (.D(branch_target_x_31__N_1122[9]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[11])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i11.GSR = "ENABLED";
    LUT4 i2_2_lut_3_lut_adj_303 (.A(csr_x[2]), .B(csr_x[1]), .C(eba[10]), 
         .Z(n3_adj_3804)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut_adj_303.init = 16'h8080;
    LUT4 i2_2_lut_3_lut_adj_304 (.A(csr_x[2]), .B(csr_x[1]), .C(eba[30]), 
         .Z(n3_adj_3805)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut_adj_304.init = 16'h8080;
    LUT4 write_idx_w_4__I_0_i3_2_lut (.A(n42732), .B(read_idx_1_d[2]), .Z(n3_adj_3806)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1490[18:47])
    defparam write_idx_w_4__I_0_i3_2_lut.init = 16'h6666;
    LUT4 i2_2_lut_3_lut_adj_305 (.A(csr_x[2]), .B(csr_x[1]), .C(eba[12]), 
         .Z(n3_adj_3807)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut_adj_305.init = 16'h8080;
    LUT4 i2_2_lut_3_lut_adj_306 (.A(csr_x[2]), .B(csr_x[1]), .C(eba[23]), 
         .Z(n3_adj_3808)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut_adj_306.init = 16'h8080;
    LUT4 i2_2_lut_3_lut_adj_307 (.A(csr_x[2]), .B(csr_x[1]), .C(eba[16]), 
         .Z(n3_adj_3809)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut_adj_307.init = 16'h8080;
    LUT4 i2_2_lut_3_lut_adj_308 (.A(csr_x[2]), .B(csr_x[1]), .C(eba[19]), 
         .Z(n3_adj_3810)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut_adj_308.init = 16'h8080;
    LUT4 mux_389_i29_3_lut (.A(branch_target_d[30]), .B(bypass_data_0[30]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i29_3_lut.init = 16'hcaca;
    LUT4 mux_389_i28_3_lut (.A(branch_target_d[29]), .B(bypass_data_0[29]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i28_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_3_lut_adj_309 (.A(csr_x[2]), .B(csr_x[1]), .C(eba[15]), 
         .Z(n3_adj_3811)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut_adj_309.init = 16'h8080;
    LUT4 i2_2_lut_3_lut_adj_310 (.A(csr_x[2]), .B(csr_x[1]), .C(eba[9]), 
         .Z(n3_adj_3812)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut_adj_310.init = 16'h8080;
    LUT4 i2_2_lut_3_lut_adj_311 (.A(csr_x[2]), .B(csr_x[1]), .C(eba[18]), 
         .Z(n3_adj_3813)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut_adj_311.init = 16'h8080;
    LUT4 i2_2_lut_3_lut_adj_312 (.A(csr_x[2]), .B(csr_x[1]), .C(eba[14]), 
         .Z(n3_adj_3814)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut_adj_312.init = 16'h8080;
    LUT4 i2_2_lut_3_lut_adj_313 (.A(csr_x[2]), .B(csr_x[1]), .C(eba[25]), 
         .Z(n3_adj_3815)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut_adj_313.init = 16'h8080;
    LUT4 mux_75_i30_3_lut (.A(logic_result_x[29]), .B(mc_result_x[29]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i30_3_lut.init = 16'hcaca;
    LUT4 mux_20532_i19_3_lut (.A(n23070), .B(n23102), .C(read_idx_0_d[4]), 
         .Z(n23116[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i19_3_lut.init = 16'hcaca;
    LUT4 mux_20532_i20_3_lut (.A(n23071), .B(n23103), .C(read_idx_0_d[4]), 
         .Z(n23116[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i20_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_3_lut_adj_314 (.A(csr_x[2]), .B(csr_x[1]), .C(eba[26]), 
         .Z(n3_adj_3776)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut_adj_314.init = 16'h8080;
    LUT4 i2_2_lut_3_lut_adj_315 (.A(csr_x[2]), .B(csr_x[1]), .C(eba[29]), 
         .Z(n3)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut_adj_315.init = 16'h8080;
    LUT4 mux_76_i18_3_lut (.A(n1253[17]), .B(sext_result_x[15]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i18_3_lut.init = 16'hcaca;
    LUT4 m_result_31__I_0_i9_3_lut (.A(m_result[8]), .B(operand_w_31__N_1187[8]), 
         .C(n42746), .Z(operand_w_31__N_840[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 mux_76_i17_3_lut (.A(n1253[16]), .B(sext_result_x[15]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i17_3_lut.init = 16'hcaca;
    LUT4 i2_2_lut_3_lut_adj_316 (.A(csr_x[2]), .B(csr_x[1]), .C(eba[31]), 
         .Z(n3_adj_3816)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i2_2_lut_3_lut_adj_316.init = 16'h8080;
    LUT4 mux_19174_i7_3_lut (.A(pc_m[8]), .B(memop_pc_w[8]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i7_3_lut.init = 16'hcaca;
    LUT4 mux_20532_i21_3_lut (.A(n23072), .B(n23104), .C(read_idx_0_d[4]), 
         .Z(n23116[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i21_3_lut.init = 16'hcaca;
    LUT4 write_enable_w_I_0_2_lut_rep_444 (.A(write_enable_w), .B(valid_w), 
         .Z(n41531)) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2015[27:74])
    defparam write_enable_w_I_0_2_lut_rep_444.init = 16'h8888;
    LUT4 mux_465_i8_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[9]), .C(eba[9]), 
         .Z(n41544)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i8_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 i20528_2_lut_rep_383_3_lut (.A(write_enable_w), .B(valid_w), .C(\counter[2] ), 
         .Z(n41470)) /* synthesis lut_function=(A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2015[27:74])
    defparam i20528_2_lut_rep_383_3_lut.init = 16'h8080;
    LUT4 i20572_2_lut_3_lut_4_lut (.A(write_enable_w), .B(valid_w), .C(write_idx_w[4]), 
         .D(\counter[2] ), .Z(n23185)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2015[27:74])
    defparam i20572_2_lut_3_lut_4_lut.init = 16'h0800;
    LUT4 mux_76_i16_3_lut (.A(n1253[15]), .B(sext_result_x[15]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i16_3_lut.init = 16'hcaca;
    LUT4 i20573_2_lut_3_lut_4_lut (.A(write_enable_w), .B(valid_w), .C(write_idx_w[4]), 
         .D(\counter[2] ), .Z(n23186)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2015[27:74])
    defparam i20573_2_lut_3_lut_4_lut.init = 16'h8000;
    PFUMX i38591 (.BLUT(n41570), .ALUT(n41571), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[15]));
    LUT4 mux_465_i8_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[9]), .C(branch_target_x[9]), 
         .Z(n41543)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i8_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    CCU2D pc_d_31__I_0_30 (.A0(pc_d[30]), .B0(instruction_d[31]), .C0(read_idx_0_d[4]), 
          .D0(instruction_d[15]), .A1(pc_d[31]), .B1(instruction_d[31]), 
          .C1(read_idx_0_d[4]), .D1(instruction_d[15]), .CIN(n36634), 
          .S0(branch_target_d[30]), .S1(branch_target_d[31]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam pc_d_31__I_0_30.INIT0 = 16'h596a;
    defparam pc_d_31__I_0_30.INIT1 = 16'h596a;
    defparam pc_d_31__I_0_30.INJECT1_0 = "NO";
    defparam pc_d_31__I_0_30.INJECT1_1 = "NO";
    FD1P3AX valid_f_617 (.D(n42726), .SP(valid_f_N_1227), .CK(w_clk_cpu), 
            .Q(valid_f)) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2264[5] 2299[8])
    defparam valid_f_617.GSR = "ENABLED";
    FD1P3AX valid_m_620 (.D(n23901), .SP(w_clk_cpu_enable_972), .CK(w_clk_cpu), 
            .Q(valid_m)) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2264[5] 2299[8])
    defparam valid_m_620.GSR = "ENABLED";
    LUT4 i36579_4_lut (.A(write_idx_w[1]), .B(write_idx_w[4]), .C(read_idx_1_d[1]), 
         .D(read_idx_1_d[4]), .Z(n39126)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i36579_4_lut.init = 16'h7bde;
    FD1P3AX store_operand_x_i0_i0 (.D(bypass_data_1[0]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[0])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i0.GSR = "ENABLED";
    FD1P3AX branch_target_x_i2_i2 (.D(branch_target_x_31__N_1122[0]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[2])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i2.GSR = "ENABLED";
    PFUMX w_result_31__I_0_i13 (.BLUT(w_result_31__N_680[12]), .ALUT(load_data_w[12]), 
          .C0(w_result_sel_load_w), .Z(w_result[12])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX csr_x_i0_i0 (.D(read_idx_0_d[0]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(csr_x[0])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam csr_x_i0_i0.GSR = "ENABLED";
    FD1P3AX eba_i8_i8 (.D(operand_1_x[8]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[8])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i8.GSR = "ENABLED";
    LUT4 mux_20532_i22_3_lut (.A(n23073), .B(n23105), .C(read_idx_0_d[4]), 
         .Z(n23116[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i22_3_lut.init = 16'hcaca;
    LUT4 mux_76_i8_3_lut (.A(n1253[7]), .B(muliplicand[7]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i8_3_lut.init = 16'hcaca;
    LUT4 mux_20532_i23_3_lut (.A(n23074), .B(n23106), .C(read_idx_0_d[4]), 
         .Z(n23116[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i23_3_lut.init = 16'hcaca;
    CCU2D pc_d_31__I_0_28 (.A0(pc_d[28]), .B0(instruction_d[31]), .C0(read_idx_0_d[4]), 
          .D0(instruction_d[15]), .A1(pc_d[29]), .B1(instruction_d[31]), 
          .C1(read_idx_0_d[4]), .D1(instruction_d[15]), .CIN(n36633), 
          .COUT(n36634), .S0(branch_target_d[28]), .S1(branch_target_d[29]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam pc_d_31__I_0_28.INIT0 = 16'h596a;
    defparam pc_d_31__I_0_28.INIT1 = 16'h596a;
    defparam pc_d_31__I_0_28.INJECT1_0 = "NO";
    defparam pc_d_31__I_0_28.INJECT1_1 = "NO";
    LUT4 mux_465_i9_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[10]), .C(eba[10]), 
         .Z(n41547)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i9_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 m_result_31__I_0_i8_3_lut (.A(m_result[7]), .B(operand_w_31__N_1187[7]), 
         .C(n42746), .Z(operand_w_31__N_840[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 mux_19174_i6_3_lut (.A(pc_m[7]), .B(memop_pc_w[7]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i6_3_lut.init = 16'hcaca;
    LUT4 mux_76_i7_3_lut (.A(n1253[6]), .B(muliplicand[6]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i7_3_lut.init = 16'hcaca;
    FD1S3IX operand_w_i0 (.D(m_result[0]), .CK(w_clk_cpu), .CD(exception_m), 
            .Q(operand_w[0])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i0.GSR = "ENABLED";
    LUT4 mux_389_i27_3_lut (.A(branch_target_d[28]), .B(bypass_data_0[28]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i27_3_lut.init = 16'hcaca;
    LUT4 mux_389_i26_3_lut (.A(branch_target_d[27]), .B(bypass_data_0[27]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i26_3_lut.init = 16'hcaca;
    LUT4 mux_76_i6_3_lut (.A(n1253[5]), .B(muliplicand[5]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i6_3_lut.init = 16'hcaca;
    FD1S3AX write_idx_w_i0 (.D(write_idx_m[0]), .CK(w_clk_cpu), .Q(write_idx_w[0])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_w_i0.GSR = "ENABLED";
    FD1S3AX w_result_sel_load_w_678 (.D(w_result_sel_load_m), .CK(w_clk_cpu), 
            .Q(w_result_sel_load_w)) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam w_result_sel_load_w_678.GSR = "ENABLED";
    FD1S3AX w_result_sel_mul_w_679 (.D(w_result_sel_mul_m), .CK(w_clk_cpu), 
            .Q(w_result_sel_mul_w)) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam w_result_sel_mul_w_679.GSR = "ENABLED";
    FD1P3AX deba_i8_i8 (.D(operand_1_x[8]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[8])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i8.GSR = "ENABLED";
    FD1S3AX write_enable_w_681 (.D(write_enable_m), .CK(w_clk_cpu), .Q(write_enable_w)) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_enable_w_681.GSR = "ENABLED";
    FD1S3AX debug_exception_w_682 (.D(debug_exception_m), .CK(w_clk_cpu), 
            .Q(debug_exception_w)) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam debug_exception_w_682.GSR = "ENABLED";
    FD1S3AX non_debug_exception_w_683 (.D(non_debug_exception_m), .CK(w_clk_cpu), 
            .Q(non_debug_exception_w)) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam non_debug_exception_w_683.GSR = "ENABLED";
    LUT4 mux_76_i5_3_lut (.A(n1253[4]), .B(muliplicand[4]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i5_3_lut.init = 16'hcaca;
    PFUMX i23_adj_317 (.BLUT(n3_adj_3811), .ALUT(n7_adj_3787), .C0(csr_x[3]), 
          .Z(n10_adj_3817));
    CCU2D pc_d_31__I_0_26 (.A0(pc_d[26]), .B0(instruction_d[31]), .C0(read_idx_0_d[3]), 
          .D0(instruction_d[15]), .A1(pc_d[27]), .B1(instruction_d[31]), 
          .C1(read_idx_0_d[4]), .D1(instruction_d[15]), .CIN(n36632), 
          .COUT(n36633), .S0(branch_target_d[26]), .S1(branch_target_d[27]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam pc_d_31__I_0_26.INIT0 = 16'h596a;
    defparam pc_d_31__I_0_26.INIT1 = 16'h596a;
    defparam pc_d_31__I_0_26.INJECT1_0 = "NO";
    defparam pc_d_31__I_0_26.INJECT1_1 = "NO";
    PFUMX w_result_31__I_0_i14 (.BLUT(w_result_31__N_680[13]), .ALUT(load_data_w[13]), 
          .C0(w_result_sel_load_w), .Z(w_result[13])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_76_i1_3_lut (.A(n1253[0]), .B(muliplicand[0]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i1_3_lut.init = 16'hcaca;
    PFUMX i38589 (.BLUT(n41567), .ALUT(n41568), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[14]));
    LUT4 x_result_31__I_17_i15_3_lut (.A(x_result_31__N_1066[14]), .B(adder_result_x[14]), 
         .C(x_result_sel_add_x), .Z(x_result_31__N_616[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam x_result_31__I_17_i15_3_lut.init = 16'hcaca;
    PFUMX w_result_31__I_0_i15 (.BLUT(w_result_31__N_680[14]), .ALUT(load_data_w[14]), 
          .C0(w_result_sel_load_w), .Z(w_result[14])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX branch_target_x_i2_i10 (.D(branch_target_x_31__N_1122[8]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[10])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i10.GSR = "ENABLED";
    FD1P3AX branch_target_x_i2_i9 (.D(branch_target_x_31__N_1122[7]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[9])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i9.GSR = "ENABLED";
    LUT4 m_result_31__I_0_i7_3_lut (.A(m_result[6]), .B(operand_w_31__N_1187[6]), 
         .C(n42746), .Z(operand_w_31__N_840[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 mux_19174_i5_3_lut (.A(pc_m[6]), .B(memop_pc_w[6]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i5_3_lut.init = 16'hcaca;
    LUT4 x_result_31__I_17_i14_3_lut (.A(x_result_31__N_1066[13]), .B(adder_result_x[13]), 
         .C(x_result_sel_add_x), .Z(x_result_31__N_616[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam x_result_31__I_17_i14_3_lut.init = 16'hcaca;
    LUT4 mux_20532_i24_3_lut (.A(n23075), .B(n23107), .C(read_idx_0_d[4]), 
         .Z(n23116[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i24_3_lut.init = 16'hcaca;
    PFUMX i23_adj_318 (.BLUT(n3_adj_3810), .ALUT(n7_adj_3786), .C0(csr_x[3]), 
          .Z(n10_adj_3818));
    LUT4 mux_20532_i25_3_lut (.A(n23076), .B(n23108), .C(read_idx_0_d[4]), 
         .Z(n23116[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i25_3_lut.init = 16'hcaca;
    LUT4 m_result_31__I_0_i6_3_lut (.A(m_result[5]), .B(operand_w_31__N_1187[5]), 
         .C(n42746), .Z(operand_w_31__N_840[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i6_3_lut.init = 16'hcaca;
    LUT4 mux_19174_i4_3_lut (.A(pc_m[5]), .B(memop_pc_w[5]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i4_3_lut.init = 16'hcaca;
    LUT4 x_result_31__I_17_i13_3_lut (.A(x_result_31__N_1066[12]), .B(adder_result_x[12]), 
         .C(x_result_sel_add_x), .Z(x_result_31__N_616[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam x_result_31__I_17_i13_3_lut.init = 16'hcaca;
    LUT4 mux_75_i25_3_lut (.A(logic_result_x[24]), .B(mc_result_x[24]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i25_3_lut.init = 16'hcaca;
    LUT4 x_result_31__I_17_i12_3_lut (.A(x_result_31__N_1066[11]), .B(adder_result_x[11]), 
         .C(x_result_sel_add_x), .Z(x_result_31__N_616[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam x_result_31__I_17_i12_3_lut.init = 16'hcaca;
    LUT4 m_result_31__I_0_i5_3_lut (.A(m_result[4]), .B(operand_w_31__N_1187[4]), 
         .C(n42746), .Z(operand_w_31__N_840[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i5_3_lut.init = 16'hcaca;
    FD1P3AX m_result_sel_compare_x_631 (.D(n41419), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(m_result_sel_compare_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam m_result_sel_compare_x_631.GSR = "ENABLED";
    LUT4 mux_19174_i3_3_lut (.A(pc_m[4]), .B(memop_pc_w[4]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i3_3_lut.init = 16'hcaca;
    PFUMX w_result_31__I_0_i16 (.BLUT(w_result_31__N_680[15]), .ALUT(load_data_w[15]), 
          .C0(w_result_sel_load_w), .Z(w_result[15])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 x_result_31__I_17_i11_3_lut (.A(x_result_31__N_1066[10]), .B(adder_result_x[10]), 
         .C(x_result_sel_add_x), .Z(x_result_31__N_616[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam x_result_31__I_17_i11_3_lut.init = 16'hcaca;
    FD1P3AX operand_1_x_i0_i31 (.D(d_result_1[31]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[31])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i31.GSR = "ENABLED";
    PFUMX i23_adj_319 (.BLUT(n3_adj_3808), .ALUT(n7_adj_3785), .C0(csr_x[3]), 
          .Z(n10_adj_3819));
    LUT4 x_result_31__I_17_i10_3_lut (.A(x_result_31__N_1066[9]), .B(adder_result_x[9]), 
         .C(x_result_sel_add_x), .Z(x_result_31__N_616[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam x_result_31__I_17_i10_3_lut.init = 16'hcaca;
    FD1P3AX operand_1_x_i0_i30 (.D(d_result_1[30]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[30])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i30.GSR = "ENABLED";
    FD1P3AX operand_1_x_i0_i29 (.D(d_result_1[29]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[29])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i29.GSR = "ENABLED";
    FD1P3AX operand_1_x_i0_i28 (.D(d_result_1[28]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[28])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i28.GSR = "ENABLED";
    FD1P3IX branch_target_m_i2_i4 (.D(branch_target_x[4]), .SP(w_clk_cpu_enable_985), 
            .CD(n22503), .CK(w_clk_cpu), .Q(branch_target_m[4])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i4.GSR = "ENABLED";
    LUT4 x_result_31__I_17_i9_3_lut (.A(x_result_31__N_1066[8]), .B(adder_result_x[8]), 
         .C(x_result_sel_add_x), .Z(x_result_31__N_616[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1608[18] 1621[32])
    defparam x_result_31__I_17_i9_3_lut.init = 16'hcaca;
    FD1P3AX operand_1_x_i0_i27 (.D(d_result_1[27]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[27])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i27.GSR = "ENABLED";
    PFUMX w_result_31__I_0_i17 (.BLUT(w_result_31__N_680[16]), .ALUT(load_data_w[16]), 
          .C0(w_result_sel_load_w), .Z(w_result[16])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i18 (.BLUT(w_result_31__N_680[17]), .ALUT(load_data_w[17]), 
          .C0(w_result_sel_load_w), .Z(w_result[17])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 stall_m_N_1109_I_0_4_lut (.A(n41428), .B(n42746), .C(n41147), 
         .D(n38972), .Z(branch_taken_m)) /* synthesis lut_function=(!(A+!(B+(C (D))))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1655[30] 1668[31])
    defparam stall_m_N_1109_I_0_4_lut.init = 16'h5444;
    LUT4 i1_2_lut_4_lut (.A(n41530), .B(csr_x[3]), .C(csr_x[4]), .D(csr_x[0]), 
         .Z(n25563)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i1_2_lut_4_lut.init = 16'h0800;
    PFUMX i38587 (.BLUT(n41564), .ALUT(n41565), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[13]));
    LUT4 mux_76_i4_3_lut (.A(n1253[3]), .B(muliplicand[3]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i4_3_lut.init = 16'hcaca;
    PFUMX w_result_31__I_0_i19 (.BLUT(w_result_31__N_680[18]), .ALUT(load_data_w[18]), 
          .C0(w_result_sel_load_w), .Z(w_result[18])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    CCU2D pc_d_31__I_0_24 (.A0(pc_d[24]), .B0(instruction_d[31]), .C0(read_idx_0_d[1]), 
          .D0(instruction_d[15]), .A1(pc_d[25]), .B1(instruction_d[31]), 
          .C1(read_idx_0_d[2]), .D1(instruction_d[15]), .CIN(n36631), 
          .COUT(n36632), .S0(branch_target_d[24]), .S1(branch_target_d[25]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam pc_d_31__I_0_24.INIT0 = 16'h596a;
    defparam pc_d_31__I_0_24.INIT1 = 16'h596a;
    defparam pc_d_31__I_0_24.INJECT1_0 = "NO";
    defparam pc_d_31__I_0_24.INJECT1_1 = "NO";
    PFUMX w_result_31__I_0_i20 (.BLUT(w_result_31__N_680[19]), .ALUT(load_data_w[19]), 
          .C0(w_result_sel_load_w), .Z(w_result[19])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3IX write_idx_x_i0_i1 (.D(write_idx_4__N_1770[1]), .SP(w_clk_cpu_enable_984), 
            .CD(n26142), .CK(w_clk_cpu), .Q(write_idx_x[1])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_x_i0_i1.GSR = "ENABLED";
    PFUMX w_result_31__I_0_i21 (.BLUT(w_result_31__N_680[20]), .ALUT(load_data_w[20]), 
          .C0(w_result_sel_load_w), .Z(w_result[20])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i22 (.BLUT(w_result_31__N_680[21]), .ALUT(load_data_w[21]), 
          .C0(w_result_sel_load_w), .Z(w_result[21])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX operand_1_x_i0_i26 (.D(d_result_1[26]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[26])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i26.GSR = "ENABLED";
    FD1P3AX operand_1_x_i0_i25 (.D(d_result_1[25]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[25])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i25.GSR = "ENABLED";
    FD1P3AX operand_1_x_i0_i24 (.D(d_result_1[24]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[24])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i24.GSR = "ENABLED";
    FD1P3AX operand_1_x_i0_i23 (.D(d_result_1[23]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[23])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i23.GSR = "ENABLED";
    PFUMX w_result_31__I_0_i23 (.BLUT(w_result_31__N_680[22]), .ALUT(load_data_w[22]), 
          .C0(w_result_sel_load_w), .Z(w_result[22])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX operand_1_x_i0_i22 (.D(d_result_1[22]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[22])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i22.GSR = "ENABLED";
    PFUMX w_result_31__I_0_i24 (.BLUT(w_result_31__N_680[23]), .ALUT(load_data_w[23]), 
          .C0(w_result_sel_load_w), .Z(w_result[23])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i25 (.BLUT(w_result_31__N_680[24]), .ALUT(load_data_w[24]), 
          .C0(w_result_sel_load_w), .Z(w_result[24])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i26 (.BLUT(w_result_31__N_680[25]), .ALUT(load_data_w[25]), 
          .C0(w_result_sel_load_w), .Z(w_result[25])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX operand_1_x_i0_i21 (.D(d_result_1[21]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[21])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i21.GSR = "ENABLED";
    FD1P3AX debug_exception_m_675 (.D(n41526), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(debug_exception_m));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam debug_exception_m_675.GSR = "ENABLED";
    PFUMX w_result_31__I_0_i27 (.BLUT(w_result_31__N_680[26]), .ALUT(load_data_w[26]), 
          .C0(w_result_sel_load_w), .Z(w_result[26])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 m_result_31__I_0_i4_3_lut (.A(m_result[3]), .B(operand_w_31__N_1187[3]), 
         .C(n42746), .Z(operand_w_31__N_840[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 mux_19174_i2_3_lut (.A(pc_m[3]), .B(memop_pc_w[3]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i2_3_lut.init = 16'hcaca;
    FD1P3AX m_result_sel_shift_m_662 (.D(m_result_sel_shift_x), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(m_result_sel_shift_m));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam m_result_sel_shift_m_662.GSR = "ENABLED";
    PFUMX w_result_31__I_0_i28 (.BLUT(w_result_31__N_680[27]), .ALUT(load_data_w[27]), 
          .C0(w_result_sel_load_w), .Z(w_result[27])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i29 (.BLUT(w_result_31__N_680[28]), .ALUT(load_data_w[28]), 
          .C0(w_result_sel_load_w), .Z(w_result[28])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i30 (.BLUT(w_result_31__N_680[29]), .ALUT(load_data_w[29]), 
          .C0(w_result_sel_load_w), .Z(w_result[29])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX w_result_31__I_0_i31 (.BLUT(w_result_31__N_680[30]), .ALUT(load_data_w[30]), 
          .C0(w_result_sel_load_w), .Z(w_result[30])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX i38585 (.BLUT(n41561), .ALUT(n41562), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[12]));
    FD1P3AX operand_1_x_i0_i20 (.D(d_result_1[20]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[20])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i20.GSR = "ENABLED";
    FD1P3AX operand_1_x_i0_i19 (.D(d_result_1[19]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[19])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i19.GSR = "ENABLED";
    FD1P3AX memop_pc_w_i2_i2 (.D(pc_m[2]), .SP(memop_pc_w_31__N_1219), .CK(w_clk_cpu), 
            .Q(memop_pc_w[2])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i2.GSR = "ENABLED";
    FD1P3AX operand_1_x_i0_i18 (.D(d_result_1[18]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[18])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i18.GSR = "ENABLED";
    LUT4 m_result_31__I_0_i3_3_lut (.A(m_result[2]), .B(operand_w_31__N_1187[2]), 
         .C(n42746), .Z(operand_w_31__N_840[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i3_3_lut.init = 16'hcaca;
    PFUMX w_result_31__I_0_i32 (.BLUT(w_result_31__N_680[31]), .ALUT(load_data_w[31]), 
          .C0(w_result_sel_load_w), .Z(w_result[31])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_19174_i1_3_lut (.A(pc_m[2]), .B(memop_pc_w[2]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i1_3_lut.init = 16'hcaca;
    LUT4 i21678_2_lut (.A(m_result_sel_compare_m), .B(n42746), .Z(n24298)) /* synthesis lut_function=(A+(B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam i21678_2_lut.init = 16'heeee;
    LUT4 mux_389_i25_3_lut (.A(branch_target_d[26]), .B(bypass_data_0[26]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i25_3_lut.init = 16'hcaca;
    LUT4 mux_389_i24_3_lut (.A(branch_target_d[25]), .B(bypass_data_0[25]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i24_3_lut.init = 16'hcaca;
    PFUMX d_result_sel_1_d_1__I_0_Mux_26_i3 (.BLUT(n1), .ALUT(n2), .C0(n41361), 
          .Z(d_result_1[26])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i38082_3_lut (.A(n41428), .B(branch_flushX_m_N_1116), .C(cycles_5__N_2495), 
         .Z(w_clk_cpu_enable_697)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;
    defparam i38082_3_lut.init = 16'h5454;
    LUT4 mux_75_i31_3_lut (.A(logic_result_x[30]), .B(mc_result_x[30]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i31_3_lut.init = 16'hcaca;
    PFUMX d_result_sel_1_d_1__I_0_Mux_25_i3 (.BLUT(n1_adj_3820), .ALUT(n2_adj_3821), 
          .C0(n41361), .Z(d_result_1[25])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_4_lut_adj_320 (.A(n29325), .B(im[3]), .C(n36690), .D(n38878), 
         .Z(csr_read_data_x[3])) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_adj_320.init = 16'hfefa;
    PFUMX d_result_sel_1_d_1__I_0_Mux_24_i3 (.BLUT(n1_adj_3822), .ALUT(n2_adj_3823), 
          .C0(n41361), .Z(d_result_1[24])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_389_i23_3_lut (.A(branch_target_d[24]), .B(bypass_data_0[24]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i23_3_lut.init = 16'hcaca;
    LUT4 mux_76_i9_3_lut (.A(n1253[8]), .B(csr_read_data_x[8]), .C(x_result_sel_csr_x), 
         .Z(x_result_31__N_1066[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i9_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut (.A(valid_m), .B(branch_m), .Z(n38972)) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2264[5] 2299[8])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 mux_75_i9_3_lut (.A(logic_result_x[8]), .B(mc_result_x[8]), .C(x_result_sel_mc_arith_x), 
         .Z(n1253[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i9_3_lut.init = 16'hcaca;
    LUT4 i38092_3_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .C(x_result_sel_sext_x), 
         .Z(n39497)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i38092_3_lut.init = 16'hefef;
    LUT4 bypass_data_0_31__I_15_i25_3_lut (.A(m_result[24]), .B(x_result[24]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i25_3_lut.init = 16'hcaca;
    LUT4 mux_46_i25_4_lut (.A(n23116[24]), .B(w_result[24]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[24])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i25_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_15_i24_3_lut (.A(m_result[23]), .B(x_result[23]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i24_3_lut.init = 16'hcaca;
    PFUMX d_result_sel_1_d_1__I_0_Mux_23_i3 (.BLUT(n1_adj_3824), .ALUT(n2_adj_3825), 
          .C0(n41361), .Z(d_result_1[23])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_46_i24_4_lut (.A(n23116[23]), .B(w_result[23]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[23])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i24_4_lut.init = 16'hcac0;
    LUT4 mux_389_i22_3_lut (.A(branch_target_d[23]), .B(bypass_data_0[23]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i22_3_lut.init = 16'hcaca;
    LUT4 mux_75_i32_3_lut (.A(logic_result_x[31]), .B(mc_result_x[31]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i32_3_lut.init = 16'hcaca;
    PFUMX d_result_sel_1_d_1__I_0_Mux_22_i3 (.BLUT(n1_adj_3826), .ALUT(n2_adj_3827), 
          .C0(n41361), .Z(d_result_1[22])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_76_i10_3_lut (.A(n1253[9]), .B(csr_read_data_x[9]), .C(x_result_sel_csr_x), 
         .Z(x_result_31__N_1066[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i10_3_lut.init = 16'hcaca;
    LUT4 mux_75_i10_3_lut (.A(logic_result_x[9]), .B(mc_result_x[9]), .C(x_result_sel_mc_arith_x), 
         .Z(n1253[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i10_3_lut.init = 16'hcaca;
    PFUMX d_result_sel_1_d_1__I_0_Mux_21_i3 (.BLUT(n1_adj_3828), .ALUT(n2_adj_3829), 
          .C0(n41361), .Z(d_result_1[21])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_76_i11_3_lut (.A(n1253[10]), .B(csr_read_data_x[10]), .C(x_result_sel_csr_x), 
         .Z(x_result_31__N_1066[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i11_3_lut.init = 16'hcaca;
    LUT4 mux_75_i11_3_lut (.A(logic_result_x[10]), .B(mc_result_x[10]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i11_3_lut.init = 16'hcaca;
    PFUMX d_result_sel_1_d_1__I_0_Mux_20_i3 (.BLUT(n1_adj_3830), .ALUT(n2_adj_3831), 
          .C0(n41361), .Z(d_result_1[20])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_4_lut_adj_321 (.A(im[8]), .B(csr_x[4]), .C(n38878), .D(n27), 
         .Z(csr_read_data_x[8])) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A !(B+!(D))) */ ;
    defparam i1_4_lut_adj_321.init = 16'hb3a0;
    PFUMX d_result_sel_1_d_1__I_0_Mux_19_i3 (.BLUT(n1_adj_3832), .ALUT(n2_adj_3833), 
          .C0(n41361), .Z(d_result_1[19])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_4_lut_adj_322 (.A(n26), .B(n22), .C(csr_x[3]), .D(csr_x[0]), 
         .Z(n27)) /* synthesis lut_function=(A+(B (C (D)))) */ ;
    defparam i1_4_lut_adj_322.init = 16'heaaa;
    PFUMX i23_adj_323 (.BLUT(n3_adj_3809), .ALUT(n7_adj_3784), .C0(csr_x[3]), 
          .Z(n10_adj_3834));
    LUT4 i2_4_lut_adj_324 (.A(csr_x[0]), .B(n41530), .C(n20), .D(\jtag_reg_addr_d[0] ), 
         .Z(n26)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_324.init = 16'hc4c0;
    LUT4 i45_4_lut (.A(csr_x[1]), .B(\jtag_reg_addr_d[1] ), .C(csr_x[2]), 
         .D(deba[8]), .Z(n22)) /* synthesis lut_function=(A (B (C))+!A !(C+!(D))) */ ;
    defparam i45_4_lut.init = 16'h8580;
    LUT4 i1_3_lut (.A(csr_x[3]), .B(csr_x[0]), .C(eba[8]), .Z(n20)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;
    defparam i1_3_lut.init = 16'h5151;
    LUT4 mux_465_i9_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[10]), .C(branch_target_x[10]), 
         .Z(n41546)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i9_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    PFUMX d_result_sel_1_d_1__I_0_Mux_18_i3 (.BLUT(n1_adj_3835), .ALUT(n2_adj_3836), 
          .C0(n41361), .Z(d_result_1[18])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i23454_3_lut_4_lut (.A(n41451), .B(n41372), .C(LM32D_CYC_O), 
         .D(wb_load_complete_N_2129), .Z(n26096)) /* synthesis lut_function=(!(A (C (D))+!A (B (C (D))+!B ((D)+!C)))) */ ;
    defparam i23454_3_lut_4_lut.init = 16'h0efe;
    LUT4 bypass_data_0_31__I_15_i23_3_lut (.A(m_result[22]), .B(x_result[22]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i23_3_lut.init = 16'hcaca;
    LUT4 mux_76_i12_3_lut (.A(n1253[11]), .B(csr_read_data_x[11]), .C(x_result_sel_csr_x), 
         .Z(x_result_31__N_1066[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i12_3_lut.init = 16'hcaca;
    FD1P3AX branch_target_x_i2_i8 (.D(branch_target_x_31__N_1122[6]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[8])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i8.GSR = "ENABLED";
    FD1P3AX branch_target_x_i2_i7 (.D(branch_target_x_31__N_1122[5]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[7])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i7.GSR = "ENABLED";
    LUT4 mux_75_i12_3_lut (.A(logic_result_x[11]), .B(mc_result_x[11]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i12_3_lut.init = 16'hcaca;
    FD1P3AX operand_1_x_i0_i17 (.D(d_result_1[17]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[17])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i17.GSR = "ENABLED";
    LUT4 mux_46_i23_4_lut (.A(n23116[22]), .B(w_result[22]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i23_4_lut.init = 16'hcac0;
    LUT4 mux_76_i13_3_lut (.A(n1253[12]), .B(csr_read_data_x[12]), .C(x_result_sel_csr_x), 
         .Z(x_result_31__N_1066[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i13_3_lut.init = 16'hcaca;
    LUT4 mux_75_i13_3_lut (.A(logic_result_x[12]), .B(mc_result_x[12]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i13_3_lut.init = 16'hcaca;
    LUT4 bypass_data_0_31__I_15_i22_3_lut (.A(m_result[21]), .B(x_result[21]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i22_3_lut.init = 16'hcaca;
    PFUMX d_result_sel_1_d_1__I_0_Mux_17_i3 (.BLUT(n1_adj_3837), .ALUT(n2_adj_3838), 
          .C0(n41361), .Z(d_result_1[17])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i11_3_lut_4_lut (.A(n41451), .B(n41372), .C(LM32D_CYC_O), .D(wb_load_complete_N_2129), 
         .Z(w_clk_cpu_enable_245)) /* synthesis lut_function=(A ((D)+!C)+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam i11_3_lut_4_lut.init = 16'hfe0e;
    LUT4 mux_46_i22_4_lut (.A(n23116[21]), .B(w_result[21]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i22_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_15_i21_3_lut (.A(m_result[20]), .B(x_result[20]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i21_3_lut.init = 16'hcaca;
    LUT4 mux_76_i14_3_lut (.A(n1253[13]), .B(csr_read_data_x[13]), .C(x_result_sel_csr_x), 
         .Z(x_result_31__N_1066[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i14_3_lut.init = 16'hcaca;
    LUT4 mux_75_i14_3_lut (.A(logic_result_x[13]), .B(mc_result_x[13]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i14_3_lut.init = 16'hcaca;
    FD1P3AX branch_target_x_i2_i6 (.D(branch_target_x_31__N_1122[4]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[6])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i6.GSR = "ENABLED";
    FD1P3AX branch_target_x_i2_i5 (.D(branch_target_x_31__N_1122[3]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[5])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i5.GSR = "ENABLED";
    LUT4 mux_46_i21_4_lut (.A(n23116[20]), .B(w_result[20]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i21_4_lut.init = 16'hcac0;
    FD1P3AX operand_1_x_i0_i16 (.D(d_result_1[16]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[16])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i16.GSR = "ENABLED";
    LUT4 mux_389_i21_3_lut (.A(branch_target_d[22]), .B(bypass_data_0[22]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i21_3_lut.init = 16'hcaca;
    LUT4 mux_389_i20_3_lut (.A(branch_target_d[21]), .B(bypass_data_0[21]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i20_3_lut.init = 16'hcaca;
    PFUMX d_result_sel_1_d_1__I_0_Mux_16_i3 (.BLUT(n1_adj_3839), .ALUT(n2_adj_3840), 
          .C0(n41361), .Z(d_result_1[16])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_76_i15_3_lut (.A(n1253[14]), .B(csr_read_data_x[14]), .C(x_result_sel_csr_x), 
         .Z(x_result_31__N_1066[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i15_3_lut.init = 16'hcaca;
    LUT4 mux_75_i15_3_lut (.A(logic_result_x[14]), .B(mc_result_x[14]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i15_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_325 (.A(n21231[0]), .B(n9), .C(n39068), .D(n41503), 
         .Z(csr_read_data_x[0])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_325.init = 16'hce0a;
    PFUMX d_result_sel_1_d_1__I_0_Mux_15_i3 (.BLUT(n1_adj_3841), .ALUT(n2_adj_3842), 
          .C0(n41361), .Z(d_result_1[15])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 bypass_data_0_31__I_15_i20_3_lut (.A(m_result[19]), .B(x_result[19]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i20_3_lut.init = 16'hcaca;
    LUT4 mux_46_i20_4_lut (.A(n23116[19]), .B(w_result[19]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i20_4_lut.init = 16'hcac0;
    CCU2D pc_d_31__I_0_22 (.A0(pc_d[22]), .B0(instruction_d[31]), .C0(read_idx_1_d[4]), 
          .D0(instruction_d[15]), .A1(pc_d[23]), .B1(instruction_d[31]), 
          .C1(read_idx_0_d[0]), .D1(instruction_d[15]), .CIN(n36630), 
          .COUT(n36631), .S0(branch_target_d[22]), .S1(branch_target_d[23]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam pc_d_31__I_0_22.INIT0 = 16'h596a;
    defparam pc_d_31__I_0_22.INIT1 = 16'h596a;
    defparam pc_d_31__I_0_22.INJECT1_0 = "NO";
    defparam pc_d_31__I_0_22.INJECT1_1 = "NO";
    LUT4 bypass_data_0_31__I_15_i19_3_lut (.A(m_result[18]), .B(x_result[18]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i19_3_lut.init = 16'hcaca;
    PFUMX w_result_31__I_0_i1 (.BLUT(w_result_31__N_680[0]), .ALUT(load_data_w[0]), 
          .C0(w_result_sel_load_w), .Z(w_result[0])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_3_lut_rep_324 (.A(n38764), .B(write_idx_m[1]), .C(read_idx_1_d[1]), 
         .Z(n41411)) /* synthesis lut_function=(A (B (C)+!B !(C))) */ ;
    defparam i1_3_lut_rep_324.init = 16'h8282;
    PFUMX d_result_sel_1_d_1__I_0_Mux_14_i3 (.BLUT(n1_adj_3843), .ALUT(n2_adj_3844), 
          .C0(n41361), .Z(d_result_1[14])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_4_lut_adj_326 (.A(jrx_csr_read_data[4]), .B(im[4]), .C(n25563), 
         .D(n38878), .Z(csr_read_data_x[4])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_326.init = 16'heca0;
    FD1P3AX branch_target_x_i2_i4 (.D(branch_target_x_31__N_1122[2]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[4])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i4.GSR = "ENABLED";
    FD1P3AX branch_target_x_i2_i3 (.D(branch_target_x_31__N_1122[1]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_target_x[3])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_x_i2_i3.GSR = "ENABLED";
    LUT4 i38046_2_lut_4_lut (.A(n38764), .B(write_idx_m[1]), .C(read_idx_1_d[1]), 
         .D(raw_x_1), .Z(n39329)) /* synthesis lut_function=(A (B (C+(D))+!B ((D)+!C))+!A (D)) */ ;
    defparam i38046_2_lut_4_lut.init = 16'hff82;
    LUT4 mux_46_i19_4_lut (.A(n23116[18]), .B(w_result[18]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i19_4_lut.init = 16'hcac0;
    LUT4 i1_4_lut_adj_327 (.A(im[9]), .B(n10_adj_3845), .C(n38878), .D(n4_adj_3846), 
         .Z(csr_read_data_x[9])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_327.init = 16'heca0;
    LUT4 i1_2_lut_adj_328 (.A(csr_x[4]), .B(csr_x[0]), .Z(n4_adj_3846)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_328.init = 16'h4444;
    PFUMX d_result_sel_1_d_1__I_0_Mux_13_i3 (.BLUT(n1_adj_3847), .ALUT(n2_adj_3848), 
          .C0(n41361), .Z(d_result_1[13])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 bypass_data_0_31__I_15_i18_3_lut (.A(m_result[17]), .B(x_result[17]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i18_3_lut.init = 16'hcaca;
    LUT4 mux_389_i19_3_lut (.A(branch_target_d[20]), .B(bypass_data_0[20]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i19_3_lut.init = 16'hcaca;
    LUT4 mux_389_i18_3_lut (.A(branch_target_d[19]), .B(bypass_data_0[19]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i18_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_329 (.A(im[10]), .B(n10_adj_3849), .C(n38878), .D(n4_adj_3846), 
         .Z(csr_read_data_x[10])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_329.init = 16'heca0;
    LUT4 i1_4_lut_adj_330 (.A(im[11]), .B(csr_x[4]), .C(n38878), .D(n31), 
         .Z(csr_read_data_x[11])) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A !(B+!(D))) */ ;
    defparam i1_4_lut_adj_330.init = 16'hb3a0;
    PFUMX d_result_sel_1_d_1__I_0_Mux_12_i3 (.BLUT(n1_adj_3850), .ALUT(n2_adj_3851), 
          .C0(n41361), .Z(d_result_1[12])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_4_lut_adj_331 (.A(jrx_csr_read_data[5]), .B(im[5]), .C(n25563), 
         .D(n38878), .Z(csr_read_data_x[5])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_331.init = 16'heca0;
    LUT4 mux_46_i18_4_lut (.A(n23116[17]), .B(w_result[17]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i18_4_lut.init = 16'hcac0;
    PFUMX d_result_sel_1_d_1__I_0_Mux_11_i3 (.BLUT(n1_adj_3852), .ALUT(n2_adj_3853), 
          .C0(n41361), .Z(d_result_1[11])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_4_lut_adj_332 (.A(jrx_csr_read_data[6]), .B(im[6]), .C(n25563), 
         .D(n38878), .Z(csr_read_data_x[6])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_332.init = 16'heca0;
    LUT4 i1_4_lut_adj_333 (.A(im[12]), .B(n10_adj_3854), .C(n38878), .D(n4_adj_3846), 
         .Z(csr_read_data_x[12])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_333.init = 16'heca0;
    CCU2D pc_d_31__I_0_20 (.A0(pc_d[20]), .B0(instruction_d[31]), .C0(read_idx_1_d[2]), 
          .D0(instruction_d[15]), .A1(pc_d[21]), .B1(instruction_d[31]), 
          .C1(read_idx_1_d[3]), .D1(instruction_d[15]), .CIN(n36629), 
          .COUT(n36630), .S0(branch_target_d[20]), .S1(branch_target_d[21]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam pc_d_31__I_0_20.INIT0 = 16'h596a;
    defparam pc_d_31__I_0_20.INIT1 = 16'h596a;
    defparam pc_d_31__I_0_20.INJECT1_0 = "NO";
    defparam pc_d_31__I_0_20.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_334 (.A(jrx_csr_read_data[7]), .B(im[7]), .C(n25563), 
         .D(n38878), .Z(csr_read_data_x[7])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_334.init = 16'heca0;
    LUT4 mux_75_i16_3_lut (.A(logic_result_x[15]), .B(mc_result_x[15]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i16_3_lut.init = 16'hcaca;
    LUT4 kill_f_I_0_719_2_lut_3_lut_4_lut (.A(n41375), .B(branch_taken_m), 
         .C(n39970), .D(w_clk_cpu_enable_984), .Z(valid_f_N_1227)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1690[20] 1693[45])
    defparam kill_f_I_0_719_2_lut_3_lut_4_lut.init = 16'hfeee;
    PFUMX d_result_sel_1_d_1__I_0_Mux_10_i3 (.BLUT(n1_adj_3855), .ALUT(n2_adj_3856), 
          .C0(n41361), .Z(d_result_1[10])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX i23_adj_335 (.BLUT(n3_adj_3807), .ALUT(n7_adj_3783), .C0(csr_x[3]), 
          .Z(n10_adj_3854));
    LUT4 mux_389_i17_3_lut (.A(branch_target_d[18]), .B(bypass_data_0[18]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i17_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_336 (.A(im[15]), .B(n10_adj_3817), .C(n38878), .D(n4_adj_3846), 
         .Z(csr_read_data_x[15])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_336.init = 16'heca0;
    PFUMX d_result_sel_1_d_1__I_0_Mux_9_i3 (.BLUT(n1_adj_3857), .ALUT(n2_adj_3858), 
          .C0(n41361), .Z(d_result_1[9])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_389_i16_3_lut (.A(branch_target_d[17]), .B(bypass_data_0[17]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i16_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_337 (.A(im[13]), .B(n10_adj_3859), .C(n38878), .D(n4_adj_3846), 
         .Z(csr_read_data_x[13])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_337.init = 16'heca0;
    LUT4 i1_4_lut_adj_338 (.A(im[14]), .B(n10_adj_3860), .C(n38878), .D(n4_adj_3846), 
         .Z(csr_read_data_x[14])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_338.init = 16'heca0;
    FD1P3AX scall_x_653 (.D(scall_d), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(scall_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam scall_x_653.GSR = "ENABLED";
    LUT4 mux_75_i1_3_lut (.A(logic_result_x[0]), .B(mc_result_x[0]), .C(x_result_sel_mc_arith_x), 
         .Z(n1253[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i1_3_lut.init = 16'hcaca;
    FD1P3AX deba_i8_i31 (.D(operand_1_x[31]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[31])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i31.GSR = "ENABLED";
    PFUMX d_result_sel_1_d_1__I_0_Mux_8_i3 (.BLUT(n1_adj_3861), .ALUT(n2_adj_3862), 
          .C0(n41361), .Z(d_result_1[8])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_389_i15_3_lut (.A(branch_target_d[16]), .B(bypass_data_0[16]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i15_3_lut.init = 16'hcaca;
    LUT4 bypass_data_0_31__I_15_i17_3_lut (.A(m_result[16]), .B(x_result[16]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i17_3_lut.init = 16'hcaca;
    LUT4 mux_389_i14_3_lut (.A(branch_target_d[15]), .B(bypass_data_0[15]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i14_3_lut.init = 16'hcaca;
    PFUMX d_result_sel_1_d_1__I_0_Mux_7_i3 (.BLUT(n1_adj_3863), .ALUT(n2_adj_3864), 
          .C0(n41361), .Z(d_result_1[7])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_46_i17_4_lut (.A(n23116[16]), .B(w_result[16]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i17_4_lut.init = 16'hcac0;
    FD1P3AX deba_i8_i30 (.D(operand_1_x[30]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[30])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i30.GSR = "ENABLED";
    PFUMX d_result_sel_1_d_1__I_0_Mux_6_i3 (.BLUT(n1_adj_3865), .ALUT(n2_adj_3866), 
          .C0(n41361), .Z(d_result_1[6])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_75_i17_3_lut (.A(logic_result_x[16]), .B(mc_result_x[16]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i17_3_lut.init = 16'hcaca;
    LUT4 mux_75_i2_3_lut (.A(logic_result_x[1]), .B(mc_result_x[1]), .C(x_result_sel_mc_arith_x), 
         .Z(n1253[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i2_3_lut.init = 16'hcaca;
    LUT4 mux_75_i3_3_lut (.A(logic_result_x[2]), .B(mc_result_x[2]), .C(x_result_sel_mc_arith_x), 
         .Z(n1253[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i3_3_lut.init = 16'hcaca;
    PFUMX d_result_sel_1_d_1__I_0_Mux_5_i3 (.BLUT(n1_adj_3867), .ALUT(n2_adj_3868), 
          .C0(n41361), .Z(d_result_1[5])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_4_lut_adj_339 (.A(im[16]), .B(n10_adj_3834), .C(n38878), .D(n4_adj_3846), 
         .Z(csr_read_data_x[16])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_339.init = 16'heca0;
    PFUMX d_result_sel_1_d_1__I_0_Mux_4_i3 (.BLUT(n1_adj_3869), .ALUT(n2_adj_3870), 
          .C0(n41361), .Z(d_result_1[4])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX deba_i8_i29 (.D(operand_1_x[29]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[29])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i29.GSR = "ENABLED";
    PFUMX i38581 (.BLUT(n41555), .ALUT(n41556), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[11]));
    LUT4 mux_389_i13_3_lut (.A(branch_target_d[14]), .B(bypass_data_0[14]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i13_3_lut.init = 16'hcaca;
    LUT4 mux_389_i12_3_lut (.A(branch_target_d[13]), .B(bypass_data_0[13]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i12_3_lut.init = 16'hcaca;
    FD1P3IX exception_m_669 (.D(exception_m_N_1355), .SP(w_clk_cpu_enable_972), 
            .CD(n31636), .CK(w_clk_cpu), .Q(exception_m));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam exception_m_669.GSR = "ENABLED";
    PFUMX i23_adj_340 (.BLUT(n3_adj_3805), .ALUT(n7_adj_3782), .C0(csr_x[3]), 
          .Z(n10_adj_3871));
    FD1P3AX deba_i8_i28 (.D(operand_1_x[28]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[28])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i28.GSR = "ENABLED";
    LUT4 mux_75_i4_3_lut (.A(logic_result_x[3]), .B(mc_result_x[3]), .C(x_result_sel_mc_arith_x), 
         .Z(n1253[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i4_3_lut.init = 16'hcaca;
    LUT4 mux_75_i18_3_lut (.A(logic_result_x[17]), .B(mc_result_x[17]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i18_3_lut.init = 16'hcaca;
    CCU2D pc_d_31__I_0_18 (.A0(pc_d[18]), .B0(instruction_d[31]), .C0(read_idx_1_d[0]), 
          .D0(instruction_d[15]), .A1(pc_d[19]), .B1(instruction_d[31]), 
          .C1(read_idx_1_d[1]), .D1(instruction_d[15]), .CIN(n36628), 
          .COUT(n36629), .S0(branch_target_d[18]), .S1(branch_target_d[19]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam pc_d_31__I_0_18.INIT0 = 16'h596a;
    defparam pc_d_31__I_0_18.INIT1 = 16'h596a;
    defparam pc_d_31__I_0_18.INJECT1_0 = "NO";
    defparam pc_d_31__I_0_18.INJECT1_1 = "NO";
    PFUMX d_result_sel_1_d_1__I_0_Mux_3_i3 (.BLUT(n1_adj_3872), .ALUT(n2_adj_3873), 
          .C0(n41361), .Z(d_result_1[3])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_4_lut_adj_341 (.A(im[17]), .B(csr_x[4]), .C(n38878), .D(n40567), 
         .Z(csr_read_data_x[17])) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A !(B+!(D))) */ ;
    defparam i1_4_lut_adj_341.init = 16'hb3a0;
    PFUMX d_result_sel_1_d_1__I_0_Mux_2_i3 (.BLUT(n1_adj_3874), .ALUT(n2_adj_3875), 
          .C0(n41361), .Z(d_result_1[2])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_75_i5_3_lut (.A(logic_result_x[4]), .B(mc_result_x[4]), .C(x_result_sel_mc_arith_x), 
         .Z(n1253[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i5_3_lut.init = 16'hcaca;
    PFUMX i23_adj_342 (.BLUT(n3_adj_3804), .ALUT(n7_adj_3781), .C0(csr_x[3]), 
          .Z(n10_adj_3849));
    PFUMX d_result_sel_1_d_1__I_0_Mux_1_i3 (.BLUT(n1_adj_3876), .ALUT(n2_adj_3877), 
          .C0(n41361), .Z(d_result_1[1])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX deba_i8_i27 (.D(operand_1_x[27]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[27])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i27.GSR = "ENABLED";
    PFUMX d_result_sel_1_d_1__I_0_Mux_0_i3 (.BLUT(n1_adj_3878), .ALUT(n2_adj_3879), 
          .C0(n41361), .Z(d_result_1[0])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX deba_i8_i26 (.D(operand_1_x[26]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[26])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i26.GSR = "ENABLED";
    FD1P3AX deba_i8_i25 (.D(operand_1_x[25]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[25])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i25.GSR = "ENABLED";
    LUT4 mux_75_i19_3_lut (.A(logic_result_x[18]), .B(mc_result_x[18]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i19_3_lut.init = 16'hcaca;
    LUT4 mux_389_i11_3_lut (.A(branch_target_d[12]), .B(bypass_data_0[12]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i11_3_lut.init = 16'hcaca;
    LUT4 mux_389_i10_3_lut (.A(branch_target_d[11]), .B(bypass_data_0[11]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i10_3_lut.init = 16'hcaca;
    PFUMX d_result_sel_1_d_1__I_0_Mux_31_i3 (.BLUT(n1_adj_3880), .ALUT(n36772), 
          .C0(n41361), .Z(d_result_1[31])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_75_i6_3_lut (.A(logic_result_x[5]), .B(mc_result_x[5]), .C(x_result_sel_mc_arith_x), 
         .Z(n1253[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i6_3_lut.init = 16'hcaca;
    LUT4 mux_75_i7_3_lut (.A(logic_result_x[6]), .B(mc_result_x[6]), .C(x_result_sel_mc_arith_x), 
         .Z(n1253[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i7_3_lut.init = 16'hcaca;
    LUT4 mux_75_i8_3_lut (.A(logic_result_x[7]), .B(mc_result_x[7]), .C(x_result_sel_mc_arith_x), 
         .Z(n1253[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i8_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i30_3_lut (.A(operand_w[29]), .B(multiplier_result_w[29]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i30_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_343 (.A(im[18]), .B(n10_adj_3881), .C(n38878), .D(n4_adj_3846), 
         .Z(csr_read_data_x[18])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_343.init = 16'heca0;
    PFUMX d_result_sel_1_d_1__I_0_Mux_30_i3 (.BLUT(n1_adj_3882), .ALUT(n2_adj_3883), 
          .C0(n41361), .Z(d_result_1[30])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_4_lut_adj_344 (.A(n42746), .B(condition_met_m), .C(n38972), 
         .D(n41507), .Z(branch_flushX_m_N_1116)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i1_4_lut_adj_344.init = 16'hfaea;
    LUT4 operand_w_31__I_0_i29_3_lut (.A(operand_w[28]), .B(multiplier_result_w[28]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i29_3_lut.init = 16'hcaca;
    PFUMX d_result_sel_1_d_1__I_0_Mux_29_i3 (.BLUT(n1_adj_3884), .ALUT(n2_adj_3885), 
          .C0(n41361), .Z(d_result_1[29])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_75_i20_3_lut (.A(logic_result_x[19]), .B(mc_result_x[19]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i20_3_lut.init = 16'hcaca;
    PFUMX d_result_sel_1_d_1__I_0_Mux_28_i3 (.BLUT(n1_adj_3886), .ALUT(n2_adj_3887), 
          .C0(n41361), .Z(d_result_1[28])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_4_lut_adj_345 (.A(im[19]), .B(n10_adj_3818), .C(n38878), .D(n4_adj_3846), 
         .Z(csr_read_data_x[19])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_345.init = 16'heca0;
    PFUMX d_result_sel_1_d_1__I_0_Mux_27_i3 (.BLUT(n1_adj_3888), .ALUT(n2_adj_3889), 
          .C0(n41361), .Z(d_result_1[27])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_75_i21_3_lut (.A(logic_result_x[20]), .B(mc_result_x[20]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i21_3_lut.init = 16'hcaca;
    FD1P3AX deba_i8_i24 (.D(operand_1_x[24]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[24])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i24.GSR = "ENABLED";
    LUT4 mux_465_i14_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[15]), .C(eba[15]), 
         .Z(n41565)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i14_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 i1_4_lut_adj_346 (.A(im[20]), .B(n10_adj_3890), .C(n38878), .D(n4_adj_3846), 
         .Z(csr_read_data_x[20])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_346.init = 16'heca0;
    LUT4 mux_75_i22_3_lut (.A(logic_result_x[21]), .B(mc_result_x[21]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i22_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_347 (.A(im[21]), .B(n10_adj_3891), .C(n38878), .D(n4_adj_3846), 
         .Z(csr_read_data_x[21])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_347.init = 16'heca0;
    LUT4 operand_w_31__I_0_i28_3_lut (.A(operand_w[27]), .B(multiplier_result_w[27]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i28_3_lut.init = 16'hcaca;
    FD1P3AX deba_i8_i23 (.D(operand_1_x[23]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[23])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i23.GSR = "ENABLED";
    LUT4 operand_w_31__I_0_i27_3_lut (.A(operand_w[26]), .B(multiplier_result_w[26]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i27_3_lut.init = 16'hcaca;
    PFUMX i38579 (.BLUT(n41552), .ALUT(n41553), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[10]));
    CCU2D operand_0_x_31__I_0_32 (.A0(operand_1_x[1]), .B0(muliplicand[1]), 
          .C0(operand_1_x[0]), .D0(muliplicand[0]), .A1(GND_net), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n36493), .S1(cmp_zero));
    defparam operand_0_x_31__I_0_32.INIT0 = 16'h9009;
    defparam operand_0_x_31__I_0_32.INIT1 = 16'hFFFF;
    defparam operand_0_x_31__I_0_32.INJECT1_0 = "YES";
    defparam operand_0_x_31__I_0_32.INJECT1_1 = "NO";
    LUT4 mux_75_i23_3_lut (.A(logic_result_x[22]), .B(mc_result_x[22]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i23_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i26_3_lut (.A(operand_w[25]), .B(multiplier_result_w[25]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i26_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_348 (.A(im[22]), .B(n10_adj_3802), .C(n38878), .D(n4_adj_3846), 
         .Z(csr_read_data_x[22])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_348.init = 16'heca0;
    FD1P3AX deba_i8_i22 (.D(operand_1_x[22]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[22])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i22.GSR = "ENABLED";
    LUT4 mux_75_i24_3_lut (.A(logic_result_x[23]), .B(mc_result_x[23]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i24_3_lut.init = 16'hcaca;
    FD1P3AX deba_i8_i21 (.D(operand_1_x[21]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[21])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i21.GSR = "ENABLED";
    CCU2D pc_d_31__I_0_16 (.A0(pc_d[16]), .B0(instruction_d[14]), .C0(GND_net), 
          .D0(GND_net), .A1(pc_d[17]), .B1(instruction_d[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n36627), .COUT(n36628), .S0(branch_target_d[16]), 
          .S1(branch_target_d[17]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam pc_d_31__I_0_16.INIT0 = 16'h5666;
    defparam pc_d_31__I_0_16.INIT1 = 16'h5666;
    defparam pc_d_31__I_0_16.INJECT1_0 = "NO";
    defparam pc_d_31__I_0_16.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_349 (.A(valid_x), .B(n9_adj_3892), .C(n7_adj_3893), 
         .D(n8), .Z(raw_x_1)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(472[26:38])
    defparam i1_4_lut_adj_349.init = 16'h8000;
    PFUMX bypass_data_1_31__I_0_i2 (.BLUT(bypass_data_1_31__N_1034[1]), .ALUT(bypass_data_1_31__N_904[1]), 
          .C0(n39329), .Z(bypass_data_1[1])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_4_lut_adj_350 (.A(im[23]), .B(n10_adj_3819), .C(n38878), .D(n4_adj_3846), 
         .Z(csr_read_data_x[23])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_350.init = 16'heca0;
    CCU2D pc_d_31__I_0_14 (.A0(pc_d[14]), .B0(instruction_d[12]), .C0(GND_net), 
          .D0(GND_net), .A1(pc_d[15]), .B1(instruction_d[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n36626), .COUT(n36627), .S0(branch_target_d[14]), 
          .S1(branch_target_d[15]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam pc_d_31__I_0_14.INIT0 = 16'h5666;
    defparam pc_d_31__I_0_14.INIT1 = 16'h5666;
    defparam pc_d_31__I_0_14.INJECT1_0 = "NO";
    defparam pc_d_31__I_0_14.INJECT1_1 = "NO";
    PFUMX bypass_data_1_31__I_0_i3 (.BLUT(bypass_data_1_31__N_1034[2]), .ALUT(bypass_data_1_31__N_904[2]), 
          .C0(n39329), .Z(bypass_data_1[2])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AY deba_i8_i20 (.D(operand_1_x[20]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[20])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i20.GSR = "ENABLED";
    LUT4 bypass_data_0_31__I_15_i16_3_lut (.A(m_result[15]), .B(x_result[15]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i16_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_351 (.A(im[24]), .B(n10_adj_3894), .C(n38878), .D(n4_adj_3846), 
         .Z(csr_read_data_x[24])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_351.init = 16'heca0;
    LUT4 mux_46_i16_4_lut (.A(n23116[15]), .B(w_result[15]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[15])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i16_4_lut.init = 16'hcac0;
    FD1P3AX deba_i8_i19 (.D(operand_1_x[19]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[19])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i19.GSR = "ENABLED";
    PFUMX bypass_data_1_31__I_0_i4 (.BLUT(bypass_data_1_31__N_1034[3]), .ALUT(bypass_data_1_31__N_904[3]), 
          .C0(n39329), .Z(bypass_data_1[3])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 bypass_data_0_31__I_15_i7_3_lut (.A(m_result[6]), .B(x_result[6]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i7_3_lut.init = 16'hcaca;
    LUT4 mux_46_i7_4_lut (.A(n23116[6]), .B(w_result[6]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[6])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i7_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_15_i8_3_lut (.A(m_result[7]), .B(x_result[7]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i8_3_lut.init = 16'hcaca;
    LUT4 mux_46_i8_4_lut (.A(n23116[7]), .B(w_result[7]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[7])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i8_4_lut.init = 16'hcac0;
    PFUMX i38577 (.BLUT(n41549), .ALUT(n41550), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[9]));
    PFUMX bypass_data_1_31__I_0_i5 (.BLUT(bypass_data_1_31__N_1034[4]), .ALUT(bypass_data_1_31__N_904[4]), 
          .C0(n39329), .Z(bypass_data_1[4])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i6 (.BLUT(bypass_data_1_31__N_1034[5]), .ALUT(bypass_data_1_31__N_904[5]), 
          .C0(n39329), .Z(bypass_data_1[5])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 bypass_data_0_31__I_15_i6_3_lut (.A(m_result[5]), .B(x_result[5]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i6_3_lut.init = 16'hcaca;
    FD1P3AX store_operand_x_i0_i31 (.D(bypass_data_1[31]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[31])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i31.GSR = "ENABLED";
    LUT4 mux_46_i6_4_lut (.A(n23116[5]), .B(w_result[5]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[5])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i6_4_lut.init = 16'hcac0;
    FD1P3AX deba_i8_i18 (.D(operand_1_x[18]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[18])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i18.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_352 (.A(im[25]), .B(n10_adj_3895), .C(n38878), .D(n4_adj_3846), 
         .Z(csr_read_data_x[25])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_352.init = 16'heca0;
    LUT4 i1_4_lut_adj_353 (.A(im[26]), .B(n10_adj_3778), .C(n38878), .D(n4_adj_3846), 
         .Z(csr_read_data_x[26])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_353.init = 16'heca0;
    PFUMX bypass_data_1_31__I_0_i7 (.BLUT(bypass_data_1_31__N_1034[6]), .ALUT(bypass_data_1_31__N_904[6]), 
          .C0(n39329), .Z(bypass_data_1[6])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 bypass_data_0_31__I_15_i5_3_lut (.A(m_result[4]), .B(x_result[4]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i5_3_lut.init = 16'hcaca;
    PFUMX bypass_data_1_31__I_0_i8 (.BLUT(bypass_data_1_31__N_1034[7]), .ALUT(bypass_data_1_31__N_904[7]), 
          .C0(n39329), .Z(bypass_data_1[7])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_46_i5_4_lut (.A(n23116[4]), .B(w_result[4]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i5_4_lut.init = 16'hcac0;
    PFUMX i23_adj_354 (.BLUT(n3_adj_3803), .ALUT(n7_adj_3780), .C0(csr_x[3]), 
          .Z(n10_adj_3859));
    PFUMX i23_adj_355 (.BLUT(n3_adj_3797), .ALUT(n7_adj_3795), .C0(csr_x[3]), 
          .Z(n10_adj_3890));
    FD1P3AX store_operand_x_i0_i30 (.D(bypass_data_1[30]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[30])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i30.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_356 (.A(im[27]), .B(csr_x[4]), .C(n38878), .D(n41321), 
         .Z(csr_read_data_x[27])) /* synthesis lut_function=(A (B (C)+!B (C+(D)))+!A !(B+!(D))) */ ;
    defparam i1_4_lut_adj_356.init = 16'hb3a0;
    LUT4 i1_4_lut_adj_357 (.A(im[28]), .B(n10_adj_3896), .C(n38878), .D(n4_adj_3846), 
         .Z(csr_read_data_x[28])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_357.init = 16'heca0;
    FD1P3AX store_operand_x_i0_i29 (.D(bypass_data_1[29]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[29])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i29.GSR = "ENABLED";
    FD1P3AX deba_i8_i17 (.D(operand_1_x[17]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[17])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i17.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_358 (.A(im[29]), .B(n10), .C(n38878), .D(n4_adj_3846), 
         .Z(csr_read_data_x[29])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_358.init = 16'heca0;
    FD1P3AX store_operand_x_i0_i28 (.D(bypass_data_1[28]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[28])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i28.GSR = "ENABLED";
    LUT4 operand_m_31__I_0_704_i1_3_lut (.A(operand_m[0]), .B(condition_met_m), 
         .C(m_result_sel_compare_m), .Z(m_result_31__N_648[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1629[18] 1631[27])
    defparam operand_m_31__I_0_704_i1_3_lut.init = 16'hcaca;
    LUT4 mux_76_i3_3_lut (.A(n1253[2]), .B(muliplicand[2]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i3_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i1_3_lut (.A(operand_w[0]), .B(multiplier_result_w[0]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i1_3_lut.init = 16'hcaca;
    FD1P3AX store_operand_x_i0_i27 (.D(bypass_data_1[27]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[27])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i27.GSR = "ENABLED";
    FD1P3AX deba_i8_i16 (.D(operand_1_x[16]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[16])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i16.GSR = "ENABLED";
    FD1P3AX memop_pc_w_i2_i31 (.D(pc_m[31]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[31])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i31.GSR = "ENABLED";
    LUT4 mux_76_i2_3_lut (.A(n1253[1]), .B(muliplicand[1]), .C(x_result_sel_sext_x), 
         .Z(x_result_31__N_1066[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1610[18] 1621[32])
    defparam mux_76_i2_3_lut.init = 16'hcaca;
    FD1P3AX memop_pc_w_i2_i30 (.D(pc_m[30]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[30])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i30.GSR = "ENABLED";
    FD1P3AX store_operand_x_i0_i26 (.D(bypass_data_1[26]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[26])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i26.GSR = "ENABLED";
    PFUMX i23_adj_359 (.BLUT(n3_adj_3799), .ALUT(n7_adj_3794), .C0(csr_x[3]), 
          .Z(n10_adj_3894));
    PFUMX bypass_data_1_31__I_0_i9 (.BLUT(bypass_data_1_31__N_1034[8]), .ALUT(bypass_data_1_31__N_904[8]), 
          .C0(n39329), .Z(bypass_data_1[8])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i10 (.BLUT(bypass_data_1_31__N_1034[9]), .ALUT(bypass_data_1_31__N_904[9]), 
          .C0(n39329), .Z(bypass_data_1[9])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_4_lut_adj_360 (.A(im[30]), .B(n10_adj_3871), .C(n38878), .D(n4_adj_3846), 
         .Z(csr_read_data_x[30])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_360.init = 16'heca0;
    FD1P3AX store_operand_x_i0_i25 (.D(bypass_data_1[25]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[25])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i25.GSR = "ENABLED";
    FD1P3AX deba_i8_i15 (.D(operand_1_x[15]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[15])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i15.GSR = "ENABLED";
    FD1P3AX memop_pc_w_i2_i29 (.D(pc_m[29]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[29])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i29.GSR = "ENABLED";
    FD1P3AX memop_pc_w_i2_i28 (.D(pc_m[28]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[28])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i28.GSR = "ENABLED";
    PFUMX bypass_data_1_31__I_0_i11 (.BLUT(bypass_data_1_31__N_1034[10]), 
          .ALUT(bypass_data_1_31__N_904[10]), .C0(n39329), .Z(bypass_data_1[10])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX i38170 (.BLUT(n40566), .ALUT(n40565), .C0(csr_x[2]), .Z(n40567));
    LUT4 i1_4_lut_adj_361 (.A(im[31]), .B(n10_adj_3897), .C(n38878), .D(n4_adj_3846), 
         .Z(csr_read_data_x[31])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B (D))) */ ;
    defparam i1_4_lut_adj_361.init = 16'heca0;
    LUT4 i1_4_lut_adj_362 (.A(n41531), .B(n39056), .C(n23668), .D(n39064), 
         .Z(n18863)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_362.init = 16'h0002;
    PFUMX bypass_data_1_31__I_0_i12 (.BLUT(bypass_data_1_31__N_1034[11]), 
          .ALUT(bypass_data_1_31__N_904[11]), .C0(n39329), .Z(bypass_data_1[11])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i36513_4_lut (.A(read_idx_1_d[2]), .B(read_idx_1_d[0]), .C(n42732), 
         .D(n42738), .Z(n39056)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i36513_4_lut.init = 16'h7bde;
    LUT4 i21064_2_lut (.A(read_idx_1_d[4]), .B(write_idx_w[4]), .Z(n23668)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1490[18:78])
    defparam i21064_2_lut.init = 16'h6666;
    FD1P3AX store_operand_x_i0_i24 (.D(bypass_data_1[24]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[24])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i24.GSR = "ENABLED";
    LUT4 i36521_4_lut (.A(read_idx_1_d[3]), .B(read_idx_1_d[1]), .C(n42734), 
         .D(write_idx_w[1]), .Z(n39064)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i36521_4_lut.init = 16'h7bde;
    FD1P3AX store_operand_x_i0_i23 (.D(bypass_data_1[23]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[23])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i23.GSR = "ENABLED";
    FD1P3AX deba_i8_i14 (.D(operand_1_x[14]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[14])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i14.GSR = "ENABLED";
    FD1P3AX memop_pc_w_i2_i27 (.D(pc_m[27]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[27])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i27.GSR = "ENABLED";
    FD1P3AX memop_pc_w_i2_i26 (.D(pc_m[26]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[26])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i26.GSR = "ENABLED";
    FD1P3AX branch_x_648 (.D(branch_d), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(branch_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_x_648.GSR = "ENABLED";
    LUT4 i3_4_lut (.A(write_idx_x[2]), .B(write_idx_x[0]), .C(read_idx_1_d[2]), 
         .D(read_idx_1_d[0]), .Z(n9_adj_3892)) /* synthesis lut_function=(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(472[26:38])
    defparam i3_4_lut.init = 16'h8421;
    PFUMX bypass_data_1_31__I_0_i13 (.BLUT(bypass_data_1_31__N_1034[12]), 
          .ALUT(bypass_data_1_31__N_904[12]), .C0(n39329), .Z(bypass_data_1[12])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX i23_adj_363 (.BLUT(n3_adj_3800), .ALUT(n7_adj_3793), .C0(csr_x[3]), 
          .Z(n10_adj_3896));
    PFUMX bypass_data_1_31__I_0_i14 (.BLUT(bypass_data_1_31__N_1034[13]), 
          .ALUT(bypass_data_1_31__N_904[13]), .C0(n39329), .Z(bypass_data_1[13])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX write_idx_m_i0_i0 (.D(write_idx_m_4__N_1152[0]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(write_idx_m[0])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_m_i0_i0.GSR = "ENABLED";
    FD1P3AX store_operand_x_i0_i22 (.D(bypass_data_1[22]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[22])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i22.GSR = "ENABLED";
    FD1P3AX deba_i8_i13 (.D(operand_1_x[13]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[13])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i13.GSR = "ENABLED";
    FD1P3AX deba_i8_i12 (.D(operand_1_x[12]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[12])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i12.GSR = "ENABLED";
    FD1P3AX memop_pc_w_i2_i25 (.D(pc_m[25]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[25])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i25.GSR = "ENABLED";
    FD1P3AX store_operand_x_i0_i21 (.D(bypass_data_1[21]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[21])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i21.GSR = "ENABLED";
    PFUMX bypass_data_1_31__I_0_i15 (.BLUT(bypass_data_1_31__N_1034[14]), 
          .ALUT(bypass_data_1_31__N_904[14]), .C0(n39329), .Z(bypass_data_1[14])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i16 (.BLUT(bypass_data_1_31__N_1034[15]), 
          .ALUT(bypass_data_1_31__N_904[15]), .C0(n39329), .Z(bypass_data_1[15])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i17 (.BLUT(bypass_data_1_31__N_1034[16]), 
          .ALUT(bypass_data_1_31__N_904[16]), .C0(n39329), .Z(bypass_data_1[16])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i18 (.BLUT(bypass_data_1_31__N_1034[17]), 
          .ALUT(bypass_data_1_31__N_904[17]), .C0(n39329), .Z(bypass_data_1[17])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX deba_i8_i11 (.D(operand_1_x[11]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[11])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i11.GSR = "ENABLED";
    FD1P3AX deba_i8_i10 (.D(operand_1_x[10]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[10])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i10.GSR = "ENABLED";
    FD1P3AX memop_pc_w_i2_i24 (.D(pc_m[24]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[24])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i24.GSR = "ENABLED";
    LUT4 bypass_data_0_31__I_15_i32_3_lut (.A(m_result[31]), .B(x_result[31]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i32_3_lut.init = 16'hcaca;
    FD1P3AX store_operand_x_i0_i20 (.D(bypass_data_1[20]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[20])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i20.GSR = "ENABLED";
    LUT4 mux_46_i32_4_lut (.A(n23116[31]), .B(w_result[31]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[31])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i32_4_lut.init = 16'hcac0;
    LUT4 i1_4_lut_adj_364 (.A(write_idx_x[3]), .B(write_idx_x[1]), .C(read_idx_1_d[3]), 
         .D(read_idx_1_d[1]), .Z(n7_adj_3893)) /* synthesis lut_function=(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(472[26:38])
    defparam i1_4_lut_adj_364.init = 16'h8421;
    PFUMX bypass_data_1_31__I_0_i19 (.BLUT(bypass_data_1_31__N_1034[18]), 
          .ALUT(bypass_data_1_31__N_904[18]), .C0(n39329), .Z(bypass_data_1[18])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 bypass_data_0_31__I_15_i31_3_lut (.A(m_result[30]), .B(x_result[30]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i31_3_lut.init = 16'hcaca;
    LUT4 mux_46_i31_4_lut (.A(n23116[30]), .B(w_result[30]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[30])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i31_4_lut.init = 16'hcac0;
    PFUMX bypass_data_1_31__I_0_i20 (.BLUT(bypass_data_1_31__N_1034[19]), 
          .ALUT(bypass_data_1_31__N_904[19]), .C0(n39329), .Z(bypass_data_1[19])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 bypass_data_0_31__I_15_i30_3_lut (.A(m_result[29]), .B(x_result[29]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i30_3_lut.init = 16'hcaca;
    LUT4 mux_46_i30_4_lut (.A(n23116[29]), .B(w_result[29]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[29])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i30_4_lut.init = 16'hcac0;
    LUT4 valid_d_I_0_2_lut_rep_300 (.A(valid_d), .B(branch_taken_m), .Z(n41387)) /* synthesis lut_function=(!((B)+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1969[14:54])
    defparam valid_d_I_0_2_lut_rep_300.init = 16'h2222;
    LUT4 bypass_data_0_31__I_15_i29_3_lut (.A(m_result[28]), .B(x_result[28]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i29_3_lut.init = 16'hcaca;
    FD1P3AX store_operand_x_i0_i19 (.D(bypass_data_1[19]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[19])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i19.GSR = "ENABLED";
    FD1P3AX deba_i8_i9 (.D(operand_1_x[9]), .SP(deba_31__N_1120), .CK(w_clk_cpu), 
            .Q(deba[9])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2171[5] 2178[8])
    defparam deba_i8_i9.GSR = "ENABLED";
    LUT4 modulus_d_I_0_2_lut_rep_286_3_lut (.A(valid_d), .B(branch_taken_m), 
         .C(n25722), .Z(n41373)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1969[14:54])
    defparam modulus_d_I_0_2_lut_rep_286_3_lut.init = 16'h0202;
    PFUMX bypass_data_1_31__I_0_i21 (.BLUT(bypass_data_1_31__N_1034[20]), 
          .ALUT(bypass_data_1_31__N_904[20]), .C0(n39329), .Z(bypass_data_1[20])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX memop_pc_w_i2_i23 (.D(pc_m[23]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[23])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i23.GSR = "ENABLED";
    FD1P3AX memop_pc_w_i2_i22 (.D(pc_m[22]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[22])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i22.GSR = "ENABLED";
    FD1P3AX write_idx_x_i0_i4 (.D(write_idx_d[4]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(write_idx_x[4])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_x_i0_i4.GSR = "ENABLED";
    PFUMX bypass_data_1_31__I_0_i22 (.BLUT(bypass_data_1_31__N_1034[21]), 
          .ALUT(bypass_data_1_31__N_904[21]), .C0(n39329), .Z(bypass_data_1[21])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i2_4_lut_adj_365 (.A(write_idx_x[4]), .B(write_enable_x), .C(read_idx_1_d[4]), 
         .D(n41408), .Z(n8)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((C+(D))+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(472[26:38])
    defparam i2_4_lut_adj_365.init = 16'h0084;
    PFUMX bypass_data_1_31__I_0_i23 (.BLUT(bypass_data_1_31__N_1034[22]), 
          .ALUT(bypass_data_1_31__N_904[22]), .C0(n39329), .Z(bypass_data_1[22])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i24 (.BLUT(bypass_data_1_31__N_1034[23]), 
          .ALUT(bypass_data_1_31__N_904[23]), .C0(n39329), .Z(bypass_data_1[23])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_3_lut_4_lut (.A(valid_d), .B(branch_taken_m), .C(n25722), 
         .D(n25724), .Z(n38799)) /* synthesis lut_function=((B+(C (D)))+!A) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1969[14:54])
    defparam i1_3_lut_4_lut.init = 16'hfddd;
    LUT4 mux_46_i29_4_lut (.A(n23116[28]), .B(w_result[28]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[28])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i29_4_lut.init = 16'hcac0;
    PFUMX bypass_data_1_31__I_0_i25 (.BLUT(bypass_data_1_31__N_1034[24]), 
          .ALUT(bypass_data_1_31__N_904[24]), .C0(n39329), .Z(bypass_data_1[24])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 bypass_data_0_31__I_15_i28_3_lut (.A(m_result[27]), .B(x_result[27]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i28_3_lut.init = 16'hcaca;
    FD1P3AX store_operand_x_i0_i18 (.D(bypass_data_1[18]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[18])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i18.GSR = "ENABLED";
    LUT4 mux_46_i28_4_lut (.A(n23116[27]), .B(w_result[27]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[27])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i28_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_15_i27_3_lut (.A(m_result[26]), .B(x_result[26]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i27_3_lut.init = 16'hcaca;
    FD1P3AX store_operand_x_i0_i17 (.D(bypass_data_1[17]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[17])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i17.GSR = "ENABLED";
    FD1S3AX write_idx_w_i4 (.D(write_idx_m[4]), .CK(w_clk_cpu), .Q(write_idx_w[4])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_w_i4.GSR = "ENABLED";
    FD1P3AX memop_pc_w_i2_i21 (.D(pc_m[21]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[21])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i21.GSR = "ENABLED";
    FD1P3AX memop_pc_w_i2_i20 (.D(pc_m[20]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[20])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i20.GSR = "ENABLED";
    FD1P3AX write_idx_x_i0_i3 (.D(write_idx_d[3]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(write_idx_x[3])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_x_i0_i3.GSR = "ENABLED";
    LUT4 size_x_1__I_0_703_i3_2_lut_rep_404 (.A(condition_x[0]), .B(size_x[1]), 
         .Z(n41491)) /* synthesis lut_function=(A+(B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1576[24:49])
    defparam size_x_1__I_0_703_i3_2_lut_rep_404.init = 16'heeee;
    LUT4 mux_46_i27_4_lut (.A(n23116[26]), .B(w_result[26]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[26])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i27_4_lut.init = 16'hcac0;
    PFUMX bypass_data_1_31__I_0_i26 (.BLUT(bypass_data_1_31__N_1034[25]), 
          .ALUT(bypass_data_1_31__N_904[25]), .C0(n39329), .Z(bypass_data_1[25])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_19172_i2_3_lut_4_lut (.A(condition_x[0]), .B(size_x[1]), .C(muliplicand[9]), 
         .D(muliplicand[7]), .Z(sext_result_x[9])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1576[24:49])
    defparam mux_19172_i2_3_lut_4_lut.init = 16'hf1e0;
    PFUMX bypass_data_1_31__I_0_i27 (.BLUT(bypass_data_1_31__N_1034[26]), 
          .ALUT(bypass_data_1_31__N_904[26]), .C0(n39329), .Z(bypass_data_1[26])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX store_operand_x_i0_i16 (.D(bypass_data_1[16]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[16])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i16.GSR = "ENABLED";
    LUT4 mux_19172_i4_3_lut_4_lut (.A(condition_x[0]), .B(size_x[1]), .C(muliplicand[11]), 
         .D(muliplicand[7]), .Z(sext_result_x[11])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1576[24:49])
    defparam mux_19172_i4_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19172_i1_3_lut_4_lut (.A(condition_x[0]), .B(size_x[1]), .C(muliplicand[8]), 
         .D(muliplicand[7]), .Z(sext_result_x[8])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1576[24:49])
    defparam mux_19172_i1_3_lut_4_lut.init = 16'hf1e0;
    LUT4 bypass_data_0_31__I_15_i26_3_lut (.A(m_result[25]), .B(x_result[25]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i26_3_lut.init = 16'hcaca;
    LUT4 mux_46_i26_4_lut (.A(n23116[25]), .B(w_result[25]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[25])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i26_4_lut.init = 16'hcac0;
    FD1P3AX store_operand_x_i0_i15 (.D(bypass_data_1[15]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[15])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i15.GSR = "ENABLED";
    FD1S3AX write_idx_w_i3 (.D(write_idx_m[3]), .CK(w_clk_cpu), .Q(write_idx_w[3])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_w_i3.GSR = "ENABLED";
    FD1P3AX memop_pc_w_i2_i19 (.D(pc_m[19]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[19])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i19.GSR = "ENABLED";
    FD1P3AX memop_pc_w_i2_i18 (.D(pc_m[18]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[18])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i18.GSR = "ENABLED";
    FD1P3AX write_idx_x_i0_i2 (.D(write_idx_d[2]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(write_idx_x[2])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_x_i0_i2.GSR = "ENABLED";
    LUT4 mux_19172_i8_3_lut_4_lut (.A(condition_x[0]), .B(size_x[1]), .C(muliplicand[15]), 
         .D(muliplicand[7]), .Z(sext_result_x[15])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1576[24:49])
    defparam mux_19172_i8_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX operand_m_i0_i0 (.D(x_result[0]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(operand_m[0])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i0.GSR = "ENABLED";
    LUT4 mux_19172_i5_3_lut_4_lut (.A(condition_x[0]), .B(size_x[1]), .C(muliplicand[12]), 
         .D(muliplicand[7]), .Z(sext_result_x[12])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1576[24:49])
    defparam mux_19172_i5_3_lut_4_lut.init = 16'hf1e0;
    LUT4 operand_w_31__I_0_i25_3_lut (.A(operand_w[24]), .B(multiplier_result_w[24]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i25_3_lut.init = 16'hcaca;
    LUT4 mux_19172_i6_3_lut_4_lut (.A(condition_x[0]), .B(size_x[1]), .C(muliplicand[13]), 
         .D(muliplicand[7]), .Z(sext_result_x[13])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1576[24:49])
    defparam mux_19172_i6_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19172_i3_3_lut_4_lut (.A(condition_x[0]), .B(size_x[1]), .C(muliplicand[10]), 
         .D(muliplicand[7]), .Z(sext_result_x[10])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1576[24:49])
    defparam mux_19172_i3_3_lut_4_lut.init = 16'hf1e0;
    LUT4 mux_19172_i7_3_lut_4_lut (.A(condition_x[0]), .B(size_x[1]), .C(muliplicand[14]), 
         .D(muliplicand[7]), .Z(sext_result_x[14])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1576[24:49])
    defparam mux_19172_i7_3_lut_4_lut.init = 16'hf1e0;
    PFUMX bypass_data_1_31__I_0_i28 (.BLUT(bypass_data_1_31__N_1034[27]), 
          .ALUT(bypass_data_1_31__N_904[27]), .C0(n39329), .Z(bypass_data_1[27])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_4_lut_4_lut_4_lut (.A(condition_x[0]), .B(size_x[1]), .C(adder_result_x[0]), 
         .D(adder_result_x[1]), .Z(byte_enable_x[1])) /* synthesis lut_function=(A (B (D))+!A (B+!(C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1576[24:49])
    defparam i1_4_lut_4_lut_4_lut.init = 16'hcd44;
    LUT4 i1_4_lut_4_lut_4_lut_adj_366 (.A(condition_x[0]), .B(size_x[1]), 
         .C(adder_result_x[0]), .D(adder_result_x[1]), .Z(byte_enable_x[0])) /* synthesis lut_function=(A (B (D))+!A (B+(C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1576[24:49])
    defparam i1_4_lut_4_lut_4_lut_adj_366.init = 16'hdc44;
    LUT4 D_CYC_O_I_0_1_lut_rep_405 (.A(LM32D_CYC_O), .Z(n41492)) /* synthesis lut_function=(!(A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1789[8:27])
    defparam D_CYC_O_I_0_1_lut_rep_405.init = 16'h5555;
    FD1P3AX store_operand_x_i0_i14 (.D(bypass_data_1[14]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[14])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i14.GSR = "ENABLED";
    FD1P3AX store_operand_x_i0_i13 (.D(bypass_data_1[13]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[13])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i13.GSR = "ENABLED";
    FD1S3AX write_idx_w_i2 (.D(write_idx_m[2]), .CK(w_clk_cpu), .Q(write_idx_w[2])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_w_i2.GSR = "ENABLED";
    LUT4 mux_465_i20_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[21]), .C(eba[21]), 
         .Z(n41580)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i20_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    PFUMX bypass_data_1_31__I_0_i29 (.BLUT(bypass_data_1_31__N_1034[28]), 
          .ALUT(bypass_data_1_31__N_904[28]), .C0(n39329), .Z(bypass_data_1[28])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX memop_pc_w_i2_i17 (.D(pc_m[17]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[17])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i17.GSR = "ENABLED";
    FD1P3AX memop_pc_w_i2_i16 (.D(pc_m[16]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[16])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i16.GSR = "ENABLED";
    LUT4 mux_465_i20_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[21]), .C(branch_target_x[21]), 
         .Z(n41579)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i20_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    FD1P3AX store_operand_x_i0_i12 (.D(bypass_data_1[12]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[12])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i12.GSR = "ENABLED";
    PFUMX bypass_data_1_31__I_0_i30 (.BLUT(bypass_data_1_31__N_1034[29]), 
          .ALUT(bypass_data_1_31__N_904[29]), .C0(n39329), .Z(bypass_data_1[29])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 bypass_data_0_31__I_15_i4_3_lut (.A(m_result[3]), .B(x_result[3]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i4_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_rep_406 (.A(load_m), .B(wb_select_m), .C(wb_load_complete), 
         .Z(n41493)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i1_3_lut_rep_406.init = 16'h0808;
    LUT4 operand_w_31__I_0_i24_3_lut (.A(operand_w[23]), .B(multiplier_result_w[23]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i24_3_lut.init = 16'hcaca;
    PFUMX bypass_data_1_31__I_0_i31 (.BLUT(bypass_data_1_31__N_1034[30]), 
          .ALUT(bypass_data_1_31__N_904[30]), .C0(n39329), .Z(bypass_data_1[30])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_1_31__I_0_i32 (.BLUT(bypass_data_1_31__N_1034[31]), 
          .ALUT(bypass_data_1_31__N_904[31]), .C0(n39329), .Z(bypass_data_1[31])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_465_i21_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[22]), .C(eba[22]), 
         .Z(n41583)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i21_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    PFUMX i37223 (.BLUT(n39775), .ALUT(n39776), .C0(logic_op_x[2]), .Z(condition_met_x));
    LUT4 mux_46_i4_4_lut (.A(n23116[3]), .B(w_result[3]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[3])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i4_4_lut.init = 16'hcac0;
    LUT4 mux_465_i21_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[22]), .C(branch_target_x[22]), 
         .Z(n41582)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i21_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 bypass_data_0_31__I_15_i1_3_lut (.A(m_result[0]), .B(x_result[0]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i1_3_lut.init = 16'hcaca;
    FD1P3AX store_operand_x_i0_i11 (.D(bypass_data_1[11]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[11])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i11.GSR = "ENABLED";
    FD1S3AX write_idx_w_i1 (.D(write_idx_m[1]), .CK(w_clk_cpu), .Q(write_idx_w[1])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_w_i1.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_364_4_lut (.A(load_m), .B(wb_select_m), .C(wb_load_complete), 
         .D(n41512), .Z(n41451)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i1_2_lut_rep_364_4_lut.init = 16'h0800;
    FD1P3AX memop_pc_w_i2_i15 (.D(pc_m[15]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[15])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i15.GSR = "ENABLED";
    LUT4 mux_465_i23_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[24]), .C(eba[24]), 
         .Z(n41586)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i23_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    FD1P3AX memop_pc_w_i2_i14 (.D(pc_m[14]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[14])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i14.GSR = "ENABLED";
    FD1P3AX operand_m_i0_i31 (.D(x_result[31]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(operand_m[31])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i31.GSR = "ENABLED";
    LUT4 mux_465_i23_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[24]), .C(branch_target_x[24]), 
         .Z(n41585)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i23_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    FD1P3AX logic_op_x_i0_i3 (.D(logic_op_d[3]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(logic_op_x[3])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam logic_op_x_i0_i3.GSR = "ENABLED";
    FD1P3AX store_operand_x_i0_i10 (.D(bypass_data_1[10]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[10])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i10.GSR = "ENABLED";
    PFUMX bypass_data_1_31__I_0_i1 (.BLUT(bypass_data_1_31__N_1034[0]), .ALUT(bypass_data_1_31__N_904[0]), 
          .C0(n39329), .Z(bypass_data_1[0])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_46_i1_4_lut (.A(n23116[0]), .B(w_result[0]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i1_4_lut.init = 16'hcac0;
    PFUMX bypass_data_0_31__I_14_i2 (.BLUT(bypass_data_0_31__N_1002[1]), .ALUT(bypass_data_0_31__N_872[1]), 
          .C0(n39363), .Z(bypass_data_0[1])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_465_i14_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[15]), .C(branch_target_x[15]), 
         .Z(n41564)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i14_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    PFUMX bypass_data_0_31__I_14_i3 (.BLUT(bypass_data_0_31__N_1002[2]), .ALUT(bypass_data_0_31__N_872[2]), 
          .C0(n39363), .Z(bypass_data_0[2])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 bypass_data_0_31__I_15_i15_3_lut (.A(m_result[14]), .B(x_result[14]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i15_3_lut.init = 16'hcaca;
    LUT4 mux_46_i15_4_lut (.A(n23116[14]), .B(w_result[14]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[14])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i15_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_15_i14_3_lut (.A(m_result[13]), .B(x_result[13]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i14_3_lut.init = 16'hcaca;
    LUT4 mux_389_i9_3_lut (.A(branch_target_d[10]), .B(bypass_data_0[10]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i9_3_lut.init = 16'hcaca;
    LUT4 mux_389_i8_3_lut (.A(branch_target_d[9]), .B(bypass_data_0[9]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i8_3_lut.init = 16'hcaca;
    FD1P3AX store_operand_x_i0_i9 (.D(bypass_data_1[9]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[9])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i9.GSR = "ENABLED";
    FD1S3AX operand_w_i31 (.D(operand_w_31__N_840[31]), .CK(w_clk_cpu), 
            .Q(operand_w[31])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i31.GSR = "ENABLED";
    FD1P3AX memop_pc_w_i2_i13 (.D(pc_m[13]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[13])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i13.GSR = "ENABLED";
    LUT4 mux_465_i24_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[25]), .C(eba[25]), 
         .Z(n41589)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i24_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    FD1P3AX memop_pc_w_i2_i12 (.D(pc_m[12]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[12])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i12.GSR = "ENABLED";
    FD1P3AX operand_m_i0_i30 (.D(x_result[30]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(operand_m[30])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i30.GSR = "ENABLED";
    FD1P3AX operand_m_i0_i29 (.D(x_result[29]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(operand_m[29])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i29.GSR = "ENABLED";
    FD1P3AX logic_op_x_i0_i2 (.D(instruction[28]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(logic_op_x[2])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam logic_op_x_i0_i2.GSR = "ENABLED";
    FD1P3AX store_operand_x_i0_i8 (.D(bypass_data_1[8]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[8])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i8.GSR = "ENABLED";
    PFUMX bypass_data_0_31__I_14_i9 (.BLUT(bypass_data_0_31__N_1002[8]), .ALUT(bypass_data_0_31__N_872[8]), 
          .C0(n39363), .Z(bypass_data_0[8])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_14_i10 (.BLUT(bypass_data_0_31__N_1002[9]), 
          .ALUT(bypass_data_0_31__N_872[9]), .C0(n39363), .Z(bypass_data_0[9])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_465_i24_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[25]), .C(branch_target_x[25]), 
         .Z(n41588)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i24_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 mux_46_i14_4_lut (.A(n23116[13]), .B(w_result[13]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[13])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i14_4_lut.init = 16'hcac0;
    LUT4 mux_465_i10_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[11]), .C(eba[11]), 
         .Z(n41550)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i10_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 bypass_data_0_31__I_15_i13_3_lut (.A(m_result[12]), .B(x_result[12]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i13_3_lut.init = 16'hcaca;
    LUT4 mux_46_i13_4_lut (.A(n23116[12]), .B(w_result[12]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[12])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i13_4_lut.init = 16'hcac0;
    FD1P3AX store_operand_x_i0_i7 (.D(bypass_data_1[7]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[7])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i7.GSR = "ENABLED";
    FD1S3AX operand_w_i30 (.D(operand_w_31__N_840[30]), .CK(w_clk_cpu), 
            .Q(operand_w[30])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i30.GSR = "ENABLED";
    PFUMX bypass_data_0_31__I_14_i11 (.BLUT(bypass_data_0_31__N_1002[10]), 
          .ALUT(bypass_data_0_31__N_872[10]), .C0(n39363), .Z(bypass_data_0[10])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX memop_pc_w_i2_i11 (.D(pc_m[11]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[11])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i11.GSR = "ENABLED";
    FD1P3AX memop_pc_w_i2_i10 (.D(pc_m[10]), .SP(memop_pc_w_31__N_1219), 
            .CK(w_clk_cpu), .Q(memop_pc_w[10])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i10.GSR = "ENABLED";
    FD1P3AX operand_m_i0_i28 (.D(x_result[28]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(operand_m[28])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i28.GSR = "ENABLED";
    LUT4 operand_w_31__I_0_i23_3_lut (.A(operand_w[22]), .B(multiplier_result_w[22]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i23_3_lut.init = 16'hcaca;
    FD1P3AX operand_m_i0_i27 (.D(x_result[27]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(operand_m[27])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i27.GSR = "ENABLED";
    PFUMX bypass_data_0_31__I_14_i12 (.BLUT(bypass_data_0_31__N_1002[11]), 
          .ALUT(bypass_data_0_31__N_872[11]), .C0(n39363), .Z(bypass_data_0[11])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 bypass_data_0_31__I_15_i12_3_lut (.A(m_result[11]), .B(x_result[11]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i12_3_lut.init = 16'hcaca;
    LUT4 mux_46_i12_4_lut (.A(n23116[11]), .B(w_result[11]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[11])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i12_4_lut.init = 16'hcac0;
    LUT4 bypass_data_0_31__I_15_i11_3_lut (.A(m_result[10]), .B(x_result[10]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i11_3_lut.init = 16'hcaca;
    PFUMX bypass_data_0_31__I_14_i13 (.BLUT(bypass_data_0_31__N_1002[12]), 
          .ALUT(bypass_data_0_31__N_872[12]), .C0(n39363), .Z(bypass_data_0[12])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_46_i11_4_lut (.A(n23116[10]), .B(w_result[10]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[10])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i11_4_lut.init = 16'hcac0;
    FD1P3AX condition_x_i0_i0 (.D(size_d[0]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(condition_x[0])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam condition_x_i0_i0.GSR = "ENABLED";
    LUT4 bypass_data_0_31__I_15_i10_3_lut (.A(m_result[9]), .B(x_result[9]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i10_3_lut.init = 16'hcaca;
    FD1P3AX store_operand_x_i0_i6 (.D(bypass_data_1[6]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[6])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i6.GSR = "ENABLED";
    LUT4 mux_46_i10_4_lut (.A(n23116[9]), .B(w_result[9]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[9])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i10_4_lut.init = 16'hcac0;
    FD1P3AX store_operand_x_i0_i5 (.D(bypass_data_1[5]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[5])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i5.GSR = "ENABLED";
    FD1S3AX operand_w_i29 (.D(operand_w_31__N_840[29]), .CK(w_clk_cpu), 
            .Q(operand_w[29])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i29.GSR = "ENABLED";
    FD1P3AX memop_pc_w_i2_i9 (.D(pc_m[9]), .SP(memop_pc_w_31__N_1219), .CK(w_clk_cpu), 
            .Q(memop_pc_w[9])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i9.GSR = "ENABLED";
    FD1P3AX memop_pc_w_i2_i8 (.D(pc_m[8]), .SP(memop_pc_w_31__N_1219), .CK(w_clk_cpu), 
            .Q(memop_pc_w[8])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i8.GSR = "ENABLED";
    FD1P3AX operand_m_i0_i26 (.D(x_result[26]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(operand_m[26])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i26.GSR = "ENABLED";
    LUT4 mux_465_i25_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[26]), .C(eba[26]), 
         .Z(n41592)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i25_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    FD1P3AX operand_m_i0_i25 (.D(x_result[25]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(operand_m[25])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i25.GSR = "ENABLED";
    LUT4 i2_4_lut_adj_367 (.A(n46), .B(n41512), .C(n41493), .D(LM32D_CYC_O), 
         .Z(w_clk_cpu_enable_886)) /* synthesis lut_function=(!(A ((D)+!B)+!A (((D)+!C)+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(407[6:21])
    defparam i2_4_lut_adj_367.init = 16'h00c8;
    LUT4 bypass_data_0_31__I_15_i9_3_lut (.A(m_result[8]), .B(x_result[8]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i9_3_lut.init = 16'hcaca;
    LUT4 mux_46_i9_4_lut (.A(n23116[8]), .B(w_result[8]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[8])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i9_4_lut.init = 16'hcac0;
    LUT4 mux_465_i25_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[26]), .C(branch_target_x[26]), 
         .Z(n41591)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i25_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    PFUMX bypass_data_0_31__I_14_i14 (.BLUT(bypass_data_0_31__N_1002[13]), 
          .ALUT(bypass_data_0_31__N_872[13]), .C0(n39363), .Z(bypass_data_0[13])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    CCU2D pc_d_31__I_0_12 (.A0(pc_d[12]), .B0(instruction_d[10]), .C0(GND_net), 
          .D0(GND_net), .A1(pc_d[13]), .B1(instruction_d[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n36625), .COUT(n36626), .S0(branch_target_d[12]), 
          .S1(branch_target_d[13]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam pc_d_31__I_0_12.INIT0 = 16'h5666;
    defparam pc_d_31__I_0_12.INIT1 = 16'h5666;
    defparam pc_d_31__I_0_12.INJECT1_0 = "NO";
    defparam pc_d_31__I_0_12.INJECT1_1 = "NO";
    FD1P3AX write_idx_x_i0_i0 (.D(write_idx_d[0]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(write_idx_x[0])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_x_i0_i0.GSR = "ENABLED";
    LUT4 mux_465_i26_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[27]), .C(eba[27]), 
         .Z(n41595)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i26_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    FD1P3AX store_operand_x_i0_i4 (.D(bypass_data_1[4]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[4])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i4.GSR = "ENABLED";
    FD1P3AX store_operand_x_i0_i3 (.D(bypass_data_1[3]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[3])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i3.GSR = "ENABLED";
    FD1S3AX operand_w_i28 (.D(operand_w_31__N_840[28]), .CK(w_clk_cpu), 
            .Q(operand_w[28])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i28.GSR = "ENABLED";
    PFUMX i38575 (.BLUT(n41546), .ALUT(n41547), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[8]));
    FD1P3AX memop_pc_w_i2_i7 (.D(pc_m[7]), .SP(memop_pc_w_31__N_1219), .CK(w_clk_cpu), 
            .Q(memop_pc_w[7])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i7.GSR = "ENABLED";
    LUT4 mux_465_i26_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[27]), .C(branch_target_x[27]), 
         .Z(n41594)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i26_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    FD1P3AX memop_pc_w_i2_i6 (.D(pc_m[6]), .SP(memop_pc_w_31__N_1219), .CK(w_clk_cpu), 
            .Q(memop_pc_w[6])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i6.GSR = "ENABLED";
    FD1P3AX operand_m_i0_i24 (.D(x_result[24]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(operand_m[24])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i24.GSR = "ENABLED";
    FD1P3AX operand_m_i0_i23 (.D(x_result[23]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(operand_m[23])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i23.GSR = "ENABLED";
    LUT4 mux_465_i10_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[11]), .C(branch_target_x[11]), 
         .Z(n41549)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i10_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    PFUMX bypass_data_0_31__I_14_i15 (.BLUT(bypass_data_0_31__N_1002[14]), 
          .ALUT(bypass_data_0_31__N_872[14]), .C0(n39363), .Z(bypass_data_0[14])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 bypass_data_0_31__I_15_i3_3_lut (.A(m_result[2]), .B(x_result[2]), 
         .C(raw_x_0), .Z(bypass_data_0_31__N_872[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1518[10] 1521[36])
    defparam bypass_data_0_31__I_15_i3_3_lut.init = 16'hcaca;
    LUT4 mux_46_i3_4_lut (.A(n23116[2]), .B(w_result[2]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i3_4_lut.init = 16'hcac0;
    PFUMX bypass_data_0_31__I_14_i1 (.BLUT(bypass_data_0_31__N_1002[0]), .ALUT(bypass_data_0_31__N_872[0]), 
          .C0(n39363), .Z(bypass_data_0[0])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX store_operand_x_i0_i2 (.D(bypass_data_1[2]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[2])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i2.GSR = "ENABLED";
    LUT4 mux_46_i2_4_lut (.A(n23116[1]), .B(w_result[1]), .C(raw_w_0), 
         .D(n22885), .Z(bypass_data_0_31__N_1002[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1521[9:36])
    defparam mux_46_i2_4_lut.init = 16'hcac0;
    FD1P3AX store_operand_x_i0_i1 (.D(bypass_data_1[1]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(store_operand_x[1])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_operand_x_i0_i1.GSR = "ENABLED";
    FD1S3AX operand_w_i27 (.D(operand_w_31__N_840[27]), .CK(w_clk_cpu), 
            .Q(operand_w[27])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i27.GSR = "ENABLED";
    LUT4 mux_465_i27_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[28]), .C(eba[28]), 
         .Z(n41598)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i27_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    FD1P3AX memop_pc_w_i2_i5 (.D(pc_m[5]), .SP(memop_pc_w_31__N_1219), .CK(w_clk_cpu), 
            .Q(memop_pc_w[5])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i5.GSR = "ENABLED";
    LUT4 mux_465_i27_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[28]), .C(branch_target_x[28]), 
         .Z(n41597)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i27_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    FD1P3AX memop_pc_w_i2_i4 (.D(pc_m[4]), .SP(memop_pc_w_31__N_1219), .CK(w_clk_cpu), 
            .Q(memop_pc_w[4])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i4.GSR = "ENABLED";
    FD1P3AX operand_m_i0_i22 (.D(x_result[22]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(operand_m[22])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i22.GSR = "ENABLED";
    LUT4 mux_465_i28_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[29]), .C(eba[29]), 
         .Z(n41601)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i28_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    FD1P3AX operand_m_i0_i21 (.D(x_result[21]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(operand_m[21])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i21.GSR = "ENABLED";
    LUT4 bypass_data_1_31__I_16_i1_3_lut (.A(m_result[0]), .B(x_result[0]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i1_3_lut.init = 16'hcaca;
    LUT4 mux_52_i1_3_lut (.A(reg_data_1[0]), .B(w_result[0]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i1_3_lut.init = 16'hcaca;
    PFUMX bypass_data_0_31__I_14_i4 (.BLUT(bypass_data_0_31__N_1002[3]), .ALUT(bypass_data_0_31__N_872[3]), 
          .C0(n39363), .Z(bypass_data_0[3])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_465_i28_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[29]), .C(branch_target_x[29]), 
         .Z(n41600)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i28_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 operand_w_31__I_0_i22_3_lut (.A(operand_w[21]), .B(multiplier_result_w[21]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i22_3_lut.init = 16'hcaca;
    LUT4 bypass_data_1_31__I_16_i32_3_lut (.A(m_result[31]), .B(x_result[31]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i32_3_lut.init = 16'hcaca;
    LUT4 mux_52_i32_3_lut (.A(reg_data_1[31]), .B(w_result[31]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i32_3_lut.init = 16'hcaca;
    FD1S3AX operand_w_i26 (.D(operand_w_31__N_840[26]), .CK(w_clk_cpu), 
            .Q(operand_w[26])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i26.GSR = "ENABLED";
    LUT4 mux_465_i18_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[19]), .C(eba[19]), 
         .Z(n41604)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i18_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_465_i18_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[19]), .C(branch_target_x[19]), 
         .Z(n41603)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i18_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    FD1P3AX memop_pc_w_i2_i3 (.D(pc_m[3]), .SP(memop_pc_w_31__N_1219), .CK(w_clk_cpu), 
            .Q(memop_pc_w[3])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam memop_pc_w_i2_i3.GSR = "ENABLED";
    LUT4 bypass_data_1_31__I_16_i31_3_lut (.A(m_result[30]), .B(x_result[30]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i31_3_lut.init = 16'hcaca;
    FD1P3AX operand_m_i0_i20 (.D(x_result[20]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(operand_m[20])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i20.GSR = "ENABLED";
    LUT4 mux_465_i17_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[18]), .C(eba[18]), 
         .Z(n41607)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i17_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    FD1P3AX operand_m_i0_i19 (.D(x_result[19]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(operand_m[19])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i19.GSR = "ENABLED";
    LUT4 mux_465_i17_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[18]), .C(branch_target_x[18]), 
         .Z(n41606)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i17_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 mux_465_i29_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[30]), .C(eba[30]), 
         .Z(n41610)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i29_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_52_i31_3_lut (.A(reg_data_1[30]), .B(w_result[30]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i31_3_lut.init = 16'hcaca;
    LUT4 bypass_data_1_31__I_16_i30_3_lut (.A(m_result[29]), .B(x_result[29]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i30_3_lut.init = 16'hcaca;
    LUT4 mux_52_i30_3_lut (.A(reg_data_1[29]), .B(w_result[29]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i30_3_lut.init = 16'hcaca;
    PFUMX bypass_data_0_31__I_14_i26 (.BLUT(bypass_data_0_31__N_1002[25]), 
          .ALUT(bypass_data_0_31__N_872[25]), .C0(n39363), .Z(bypass_data_0[25])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 bypass_data_1_31__I_16_i29_3_lut (.A(m_result[28]), .B(x_result[28]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i29_3_lut.init = 16'hcaca;
    LUT4 mux_52_i29_3_lut (.A(reg_data_1[28]), .B(w_result[28]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i29_3_lut.init = 16'hcaca;
    FD1S3AX operand_w_i25 (.D(operand_w_31__N_840[25]), .CK(w_clk_cpu), 
            .Q(operand_w[25])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i25.GSR = "ENABLED";
    LUT4 mux_465_i29_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[30]), .C(branch_target_x[30]), 
         .Z(n41609)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i29_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 i21356_2_lut_rep_272_3_lut_4_lut (.A(valid_x), .B(n41408), .C(n25705), 
         .D(csr_write_enable_x), .Z(n41359)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1982[14:54])
    defparam i21356_2_lut_rep_272_3_lut_4_lut.init = 16'h0200;
    LUT4 bypass_data_1_31__I_16_i28_3_lut (.A(m_result[27]), .B(x_result[27]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i28_3_lut.init = 16'hcaca;
    FD1P3AX operand_m_i0_i18 (.D(x_result[18]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(operand_m[18])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i18.GSR = "ENABLED";
    LUT4 mux_465_i22_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[23]), .C(eba[23]), 
         .Z(n41613)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i22_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    FD1P3AX operand_m_i0_i17 (.D(x_result[17]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(operand_m[17])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i17.GSR = "ENABLED";
    PFUMX bypass_data_0_31__I_14_i27 (.BLUT(bypass_data_0_31__N_1002[26]), 
          .ALUT(bypass_data_0_31__N_872[26]), .C0(n39363), .Z(bypass_data_0[26])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_52_i28_3_lut (.A(reg_data_1[27]), .B(w_result[27]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i28_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i21_3_lut (.A(operand_w[20]), .B(multiplier_result_w[20]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i21_3_lut.init = 16'hcaca;
    PFUMX bypass_data_0_31__I_14_i28 (.BLUT(bypass_data_0_31__N_1002[27]), 
          .ALUT(bypass_data_0_31__N_872[27]), .C0(n39363), .Z(bypass_data_0[27])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_14_i29 (.BLUT(bypass_data_0_31__N_1002[28]), 
          .ALUT(bypass_data_0_31__N_872[28]), .C0(n39363), .Z(bypass_data_0[28])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_3_lut_adj_368 (.A(n38764), .B(read_idx_1_d[1]), .C(write_idx_m[1]), 
         .Z(n18869)) /* synthesis lut_function=(A (B (C)+!B !(C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(472[26:38])
    defparam i1_3_lut_adj_368.init = 16'h8282;
    FD1S3AX operand_w_i24 (.D(operand_w_31__N_840[24]), .CK(w_clk_cpu), 
            .Q(operand_w[24])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i24.GSR = "ENABLED";
    LUT4 mux_465_i22_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[23]), .C(branch_target_x[23]), 
         .Z(n41612)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i22_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 bypass_data_1_31__I_16_i27_3_lut (.A(m_result[26]), .B(x_result[26]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i27_3_lut.init = 16'hcaca;
    LUT4 mux_52_i27_3_lut (.A(reg_data_1[26]), .B(w_result[26]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i27_3_lut.init = 16'hcaca;
    FD1P3AX operand_m_i0_i16 (.D(x_result[16]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(operand_m[16])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i16.GSR = "ENABLED";
    FD1P3AX operand_m_i0_i15 (.D(x_result[15]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(operand_m[15])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i15.GSR = "ENABLED";
    PFUMX bypass_data_0_31__I_14_i30 (.BLUT(bypass_data_0_31__N_1002[29]), 
          .ALUT(bypass_data_0_31__N_872[29]), .C0(n39363), .Z(bypass_data_0[29])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 operand_w_31__I_0_i20_3_lut (.A(operand_w[19]), .B(multiplier_result_w[19]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i20_3_lut.init = 16'hcaca;
    PFUMX bypass_data_0_31__I_14_i31 (.BLUT(bypass_data_0_31__N_1002[30]), 
          .ALUT(bypass_data_0_31__N_872[30]), .C0(n39363), .Z(bypass_data_0[30])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_14_i32 (.BLUT(bypass_data_0_31__N_1002[31]), 
          .ALUT(bypass_data_0_31__N_872[31]), .C0(n39363), .Z(bypass_data_0[31])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_465_i6_4_lut (.A(branch_target_x[7]), .B(eid_x_2__N_999[2]), 
         .C(n41430), .D(reset_exception), .Z(branch_target_m_31__N_1157[5])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2555[7:45])
    defparam mux_465_i6_4_lut.init = 16'h0aca;
    LUT4 bypass_data_1_31__I_16_i26_3_lut (.A(m_result[25]), .B(x_result[25]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i26_3_lut.init = 16'hcaca;
    LUT4 mux_52_i26_3_lut (.A(reg_data_1[25]), .B(w_result[25]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i26_3_lut.init = 16'hcaca;
    FD1S3AX operand_w_i23 (.D(operand_w_31__N_840[23]), .CK(w_clk_cpu), 
            .Q(operand_w[23])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i23.GSR = "ENABLED";
    LUT4 bypass_data_1_31__I_16_i25_3_lut (.A(m_result[24]), .B(x_result[24]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i25_3_lut.init = 16'hcaca;
    FD1S3AX operand_w_i22 (.D(operand_w_31__N_840[22]), .CK(w_clk_cpu), 
            .Q(operand_w[22])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i22.GSR = "ENABLED";
    LUT4 mux_52_i25_3_lut (.A(reg_data_1[24]), .B(w_result[24]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i25_3_lut.init = 16'hcaca;
    FD1P3AX operand_m_i0_i14 (.D(x_result[14]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(operand_m[14])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i14.GSR = "ENABLED";
    LUT4 operand_w_31__I_0_i19_3_lut (.A(operand_w[18]), .B(multiplier_result_w[18]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i19_3_lut.init = 16'hcaca;
    LUT4 bypass_data_1_31__I_16_i24_3_lut (.A(m_result[23]), .B(x_result[23]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i24_3_lut.init = 16'hcaca;
    LUT4 mux_52_i24_3_lut (.A(reg_data_1[23]), .B(w_result[23]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i24_3_lut.init = 16'hcaca;
    LUT4 bypass_data_1_31__I_16_i23_3_lut (.A(m_result[22]), .B(x_result[22]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i23_3_lut.init = 16'hcaca;
    LUT4 mux_52_i23_3_lut (.A(reg_data_1[22]), .B(w_result[22]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i23_3_lut.init = 16'hcaca;
    LUT4 bypass_data_1_31__I_16_i22_3_lut (.A(m_result[21]), .B(x_result[21]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i22_3_lut.init = 16'hcaca;
    LUT4 mux_52_i22_3_lut (.A(reg_data_1[21]), .B(w_result[21]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i22_3_lut.init = 16'hcaca;
    FD1S3AX operand_w_i21 (.D(operand_w_31__N_840[21]), .CK(w_clk_cpu), 
            .Q(operand_w[21])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i21.GSR = "ENABLED";
    LUT4 bypass_data_1_31__I_16_i21_3_lut (.A(m_result[20]), .B(x_result[20]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i21_3_lut.init = 16'hcaca;
    LUT4 mux_52_i21_3_lut (.A(reg_data_1[20]), .B(w_result[20]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i21_3_lut.init = 16'hcaca;
    FD1S3AX operand_w_i20 (.D(operand_w_31__N_840[20]), .CK(w_clk_cpu), 
            .Q(operand_w[20])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i20.GSR = "ENABLED";
    LUT4 bypass_data_1_31__I_16_i20_3_lut (.A(m_result[19]), .B(x_result[19]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i20_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_4_lut_adj_369 (.A(valid_x), .B(n41408), .C(store_x), 
         .D(load_x), .Z(stall_a_N_1259)) /* synthesis lut_function=(!((B+!(C+(D)))+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1982[14:54])
    defparam i1_3_lut_4_lut_adj_369.init = 16'h2220;
    FD1P3AX operand_m_i0_i13 (.D(x_result[13]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(operand_m[13])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i13.GSR = "ENABLED";
    LUT4 i29587_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[28]), 
         .D(operand_m[28]), .Z(m_result[28])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29587_4_lut_4_lut.init = 16'h5140;
    LUT4 i29588_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[27]), 
         .D(operand_m[27]), .Z(m_result[27])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29588_4_lut_4_lut.init = 16'h5140;
    FD1S3AX operand_w_i19 (.D(operand_w_31__N_840[19]), .CK(w_clk_cpu), 
            .Q(operand_w[19])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i19.GSR = "ENABLED";
    LUT4 mux_465_i5_4_lut (.A(branch_target_x[6]), .B(n23893), .C(n41430), 
         .D(n38801), .Z(branch_target_m_31__N_1157[4])) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2555[7:45])
    defparam mux_465_i5_4_lut.init = 16'h3a0a;
    LUT4 mux_52_i20_3_lut (.A(reg_data_1[19]), .B(w_result[19]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i20_3_lut.init = 16'hcaca;
    LUT4 i29598_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[26]), 
         .D(operand_m[26]), .Z(m_result[26])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29598_4_lut_4_lut.init = 16'h5140;
    LUT4 mux_465_i4_4_lut (.A(branch_target_x[5]), .B(eid_x_2__N_1098[0]), 
         .C(n41430), .D(n23893), .Z(branch_target_m_31__N_1157[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2555[7:45])
    defparam mux_465_i4_4_lut.init = 16'h0aca;
    CCU2D pc_d_31__I_0_10 (.A0(pc_d[10]), .B0(instruction_d[8]), .C0(GND_net), 
          .D0(GND_net), .A1(pc_d[11]), .B1(instruction_d[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n36624), .COUT(n36625), .S0(branch_target_d[10]), 
          .S1(branch_target_d[11]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam pc_d_31__I_0_10.INIT0 = 16'h5666;
    defparam pc_d_31__I_0_10.INIT1 = 16'h5666;
    defparam pc_d_31__I_0_10.INJECT1_0 = "NO";
    defparam pc_d_31__I_0_10.INJECT1_1 = "NO";
    LUT4 bypass_data_1_31__I_16_i19_3_lut (.A(m_result[18]), .B(x_result[18]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i19_3_lut.init = 16'hcaca;
    LUT4 mux_52_i19_3_lut (.A(reg_data_1[18]), .B(w_result[18]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i19_3_lut.init = 16'hcaca;
    LUT4 i29608_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[24]), 
         .D(operand_m[24]), .Z(m_result[24])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29608_4_lut_4_lut.init = 16'h5140;
    LUT4 i29599_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[25]), 
         .D(operand_m[25]), .Z(m_result[25])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29599_4_lut_4_lut.init = 16'h5140;
    LUT4 i29609_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[23]), 
         .D(operand_m[23]), .Z(m_result[23])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29609_4_lut_4_lut.init = 16'h5140;
    LUT4 i29616_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[22]), 
         .D(operand_m[22]), .Z(m_result[22])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29616_4_lut_4_lut.init = 16'h5140;
    LUT4 i29617_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[21]), 
         .D(operand_m[21]), .Z(m_result[21])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29617_4_lut_4_lut.init = 16'h5140;
    LUT4 i29624_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[20]), 
         .D(operand_m[20]), .Z(m_result[20])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29624_4_lut_4_lut.init = 16'h5140;
    LUT4 bypass_data_1_31__I_16_i18_3_lut (.A(m_result[17]), .B(x_result[17]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i18_3_lut.init = 16'hcaca;
    LUT4 i29625_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[19]), 
         .D(operand_m[19]), .Z(m_result[19])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29625_4_lut_4_lut.init = 16'h5140;
    LUT4 i29636_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[18]), 
         .D(operand_m[18]), .Z(m_result[18])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29636_4_lut_4_lut.init = 16'h5140;
    FD1P3AX operand_m_i0_i12 (.D(x_result[12]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(operand_m[12])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i12.GSR = "ENABLED";
    LUT4 i29572_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[29]), 
         .D(operand_m[29]), .Z(m_result[29])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29572_4_lut_4_lut.init = 16'h5140;
    FD1P3AX operand_m_i0_i11 (.D(x_result[11]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(operand_m[11])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i11.GSR = "ENABLED";
    FD1P3AX operand_1_x_i0_i15 (.D(d_result_1[15]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(operand_1_x[15])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_1_x_i0_i15.GSR = "ENABLED";
    LUT4 mux_52_i18_3_lut (.A(reg_data_1[17]), .B(w_result[17]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i18_3_lut.init = 16'hcaca;
    LUT4 i29637_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[17]), 
         .D(operand_m[17]), .Z(m_result[17])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29637_4_lut_4_lut.init = 16'h5140;
    LUT4 i29644_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[16]), 
         .D(operand_m[16]), .Z(m_result[16])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29644_4_lut_4_lut.init = 16'h5140;
    LUT4 bypass_data_1_31__I_16_i17_3_lut (.A(m_result[16]), .B(x_result[16]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i17_3_lut.init = 16'hcaca;
    LUT4 mux_52_i17_3_lut (.A(reg_data_1[16]), .B(w_result[16]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i17_3_lut.init = 16'hcaca;
    LUT4 i29571_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[30]), 
         .D(operand_m[30]), .Z(m_result[30])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29571_4_lut_4_lut.init = 16'h5140;
    LUT4 i29559_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[31]), 
         .D(operand_m[31]), .Z(m_result[31])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29559_4_lut_4_lut.init = 16'h5140;
    LUT4 i29645_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[15]), 
         .D(operand_m[15]), .Z(m_result[15])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29645_4_lut_4_lut.init = 16'h5140;
    LUT4 i29655_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[14]), 
         .D(operand_m[14]), .Z(m_result[14])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29655_4_lut_4_lut.init = 16'h5140;
    LUT4 i29656_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[13]), 
         .D(operand_m[13]), .Z(m_result[13])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29656_4_lut_4_lut.init = 16'h5140;
    LUT4 i29665_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[12]), 
         .D(operand_m[12]), .Z(m_result[12])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29665_4_lut_4_lut.init = 16'h5140;
    LUT4 i29666_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[11]), 
         .D(operand_m[11]), .Z(m_result[11])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29666_4_lut_4_lut.init = 16'h5140;
    LUT4 bypass_data_1_31__I_16_i16_3_lut (.A(m_result[15]), .B(x_result[15]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i16_3_lut.init = 16'hcaca;
    FD1S3AX operand_w_i18 (.D(operand_w_31__N_840[18]), .CK(w_clk_cpu), 
            .Q(operand_w[18])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i18.GSR = "ENABLED";
    LUT4 mux_52_i16_3_lut (.A(reg_data_1[15]), .B(w_result[15]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i16_3_lut.init = 16'hcaca;
    LUT4 i29677_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[10]), 
         .D(operand_m[10]), .Z(m_result[10])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29677_4_lut_4_lut.init = 16'h5140;
    LUT4 i29678_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[9]), 
         .D(operand_m[9]), .Z(m_result[9])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29678_4_lut_4_lut.init = 16'h5140;
    FD1P3AX operand_m_i0_i10 (.D(x_result[10]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(operand_m[10])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i10.GSR = "ENABLED";
    FD1P3AX operand_m_i0_i9 (.D(x_result[9]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(operand_m[9])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i9.GSR = "ENABLED";
    LUT4 bypass_data_1_31__I_16_i15_3_lut (.A(m_result[14]), .B(x_result[14]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i15_3_lut.init = 16'hcaca;
    CCU2D pc_d_31__I_0_8 (.A0(pc_d[8]), .B0(instruction_d[6]), .C0(GND_net), 
          .D0(GND_net), .A1(pc_d[9]), .B1(instruction_d[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n36623), .COUT(n36624), .S0(branch_target_d[8]), 
          .S1(branch_target_d[9]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam pc_d_31__I_0_8.INIT0 = 16'h5666;
    defparam pc_d_31__I_0_8.INIT1 = 16'h5666;
    defparam pc_d_31__I_0_8.INJECT1_0 = "NO";
    defparam pc_d_31__I_0_8.INJECT1_1 = "NO";
    PFUMX x_result_31__I_0_i2 (.BLUT(x_result_31__N_1066[1]), .ALUT(x_result_31__N_616[1]), 
          .C0(n39459), .Z(x_result[1])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_52_i15_3_lut (.A(reg_data_1[14]), .B(w_result[14]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i15_3_lut.init = 16'hcaca;
    LUT4 bypass_data_1_31__I_16_i14_3_lut (.A(m_result[13]), .B(x_result[13]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i14_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_370 (.A(n34433), .B(n39886), .C(n6), .D(n39890), 
         .Z(n38764)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(472[26:38])
    defparam i1_4_lut_adj_370.init = 16'h0020;
    FD1S3AX operand_w_i17 (.D(operand_w_31__N_840[17]), .CK(w_clk_cpu), 
            .Q(operand_w[17])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i17.GSR = "ENABLED";
    PFUMX x_result_31__I_0_i3 (.BLUT(x_result_31__N_1066[2]), .ALUT(x_result_31__N_616[2]), 
          .C0(n39459), .Z(x_result[2])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX operand_m_i0_i8 (.D(x_result[8]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(operand_m[8])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i8.GSR = "ENABLED";
    LUT4 i29685_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[8]), 
         .D(operand_m[8]), .Z(m_result[8])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29685_4_lut_4_lut.init = 16'h5140;
    FD1P3AX operand_m_i0_i7 (.D(x_result[7]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(operand_m[7])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i7.GSR = "ENABLED";
    FD1S3AX operand_w_i16 (.D(operand_w_31__N_840[16]), .CK(w_clk_cpu), 
            .Q(operand_w[16])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i16.GSR = "ENABLED";
    LUT4 operand_w_31__I_0_i3_3_lut (.A(operand_w[2]), .B(multiplier_result_w[2]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i3_3_lut.init = 16'hcaca;
    CCU2D operand_0_x_31__I_0_23 (.A0(operand_1_x[21]), .B0(muliplicand[21]), 
          .C0(operand_1_x[20]), .D0(muliplicand[20]), .A1(operand_1_x[19]), 
          .B1(muliplicand[19]), .C1(operand_1_x[18]), .D1(muliplicand[18]), 
          .CIN(n36488), .COUT(n36489));
    defparam operand_0_x_31__I_0_23.INIT0 = 16'h9009;
    defparam operand_0_x_31__I_0_23.INIT1 = 16'h9009;
    defparam operand_0_x_31__I_0_23.INJECT1_0 = "YES";
    defparam operand_0_x_31__I_0_23.INJECT1_1 = "YES";
    PFUMX bypass_data_0_31__I_14_i5 (.BLUT(bypass_data_0_31__N_1002[4]), .ALUT(bypass_data_0_31__N_872[4]), 
          .C0(n39363), .Z(bypass_data_0[4])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_14_i6 (.BLUT(bypass_data_0_31__N_1002[5]), .ALUT(bypass_data_0_31__N_872[5]), 
          .C0(n39363), .Z(bypass_data_0[5])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i29686_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[7]), 
         .D(operand_m[7]), .Z(m_result[7])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29686_4_lut_4_lut.init = 16'h5140;
    CCU2D operand_0_x_31__I_0_31 (.A0(operand_1_x[5]), .B0(muliplicand[5]), 
          .C0(operand_1_x[4]), .D0(muliplicand[4]), .A1(operand_1_x[3]), 
          .B1(muliplicand[3]), .C1(operand_1_x[2]), .D1(muliplicand[2]), 
          .CIN(n36492), .COUT(n36493));
    defparam operand_0_x_31__I_0_31.INIT0 = 16'h9009;
    defparam operand_0_x_31__I_0_31.INIT1 = 16'h9009;
    defparam operand_0_x_31__I_0_31.INJECT1_0 = "YES";
    defparam operand_0_x_31__I_0_31.INJECT1_1 = "YES";
    LUT4 i29693_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[6]), 
         .D(operand_m[6]), .Z(m_result[6])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29693_4_lut_4_lut.init = 16'h5140;
    LUT4 i29694_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[5]), 
         .D(operand_m[5]), .Z(m_result[5])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29694_4_lut_4_lut.init = 16'h5140;
    FD1P3AX operand_m_i0_i6 (.D(x_result[6]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(operand_m[6])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i6.GSR = "ENABLED";
    LUT4 i29702_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[4]), 
         .D(operand_m[4]), .Z(m_result[4])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29702_4_lut_4_lut.init = 16'h5140;
    LUT4 i29703_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[3]), 
         .D(operand_m[3]), .Z(m_result[3])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29703_4_lut_4_lut.init = 16'h5140;
    LUT4 i29712_4_lut_4_lut (.A(n42730), .B(n42736), .C(shifter_result_m[2]), 
         .D(operand_m[2]), .Z(m_result[2])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i29712_4_lut_4_lut.init = 16'h5140;
    FD1P3AX operand_m_i0_i5 (.D(x_result[5]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(operand_m[5])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i5.GSR = "ENABLED";
    CCU2D operand_0_x_31__I_0_21 (.A0(operand_1_x[25]), .B0(muliplicand[25]), 
          .C0(operand_1_x[24]), .D0(muliplicand[24]), .A1(operand_1_x[23]), 
          .B1(muliplicand[23]), .C1(operand_1_x[22]), .D1(muliplicand[22]), 
          .CIN(n36487), .COUT(n36488));
    defparam operand_0_x_31__I_0_21.INIT0 = 16'h9009;
    defparam operand_0_x_31__I_0_21.INIT1 = 16'h9009;
    defparam operand_0_x_31__I_0_21.INJECT1_0 = "YES";
    defparam operand_0_x_31__I_0_21.INJECT1_1 = "YES";
    PFUMX bypass_data_0_31__I_14_i8 (.BLUT(bypass_data_0_31__N_1002[7]), .ALUT(bypass_data_0_31__N_872[7]), 
          .C0(n39363), .Z(bypass_data_0[7])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    CCU2D pc_d_31__I_0_6 (.A0(pc_d[6]), .B0(instruction_d[4]), .C0(GND_net), 
          .D0(GND_net), .A1(pc_d[7]), .B1(instruction_d[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n36622), .COUT(n36623), .S0(branch_target_d[6]), 
          .S1(branch_target_d[7]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam pc_d_31__I_0_6.INIT0 = 16'h5666;
    defparam pc_d_31__I_0_6.INIT1 = 16'h5666;
    defparam pc_d_31__I_0_6.INJECT1_0 = "NO";
    defparam pc_d_31__I_0_6.INJECT1_1 = "NO";
    CCU2D pc_d_31__I_0_4 (.A0(pc_d[4]), .B0(instruction_d[2]), .C0(GND_net), 
          .D0(GND_net), .A1(pc_d[5]), .B1(instruction_d[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n36621), .COUT(n36622), .S0(branch_target_d[4]), 
          .S1(branch_target_d[5]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam pc_d_31__I_0_4.INIT0 = 16'h5666;
    defparam pc_d_31__I_0_4.INIT1 = 16'h5666;
    defparam pc_d_31__I_0_4.INJECT1_0 = "NO";
    defparam pc_d_31__I_0_4.INJECT1_1 = "NO";
    CCU2D pc_d_31__I_0_2 (.A0(pc_d[2]), .B0(instruction_d[0]), .C0(GND_net), 
          .D0(GND_net), .A1(pc_d[3]), .B1(instruction_d[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n36621), .S1(branch_target_d[3]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1547[29:51])
    defparam pc_d_31__I_0_2.INIT0 = 16'h7000;
    defparam pc_d_31__I_0_2.INIT1 = 16'h5666;
    defparam pc_d_31__I_0_2.INJECT1_0 = "NO";
    defparam pc_d_31__I_0_2.INJECT1_1 = "NO";
    PFUMX bypass_data_0_31__I_14_i7 (.BLUT(bypass_data_0_31__N_1002[6]), .ALUT(bypass_data_0_31__N_872[6]), 
          .C0(n39363), .Z(bypass_data_0[6])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 bypass_data_1_31__I_16_i2_3_lut_4_lut_4_lut (.A(m_result_sel_compare_m), 
         .B(x_result[1]), .C(raw_x_1), .D(n41438), .Z(bypass_data_1_31__N_904[1])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam bypass_data_1_31__I_16_i2_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 mux_52_i14_3_lut (.A(reg_data_1[13]), .B(w_result[13]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i14_3_lut.init = 16'hcaca;
    LUT4 bypass_data_0_31__I_15_i2_3_lut_4_lut_4_lut (.A(m_result_sel_compare_m), 
         .B(x_result[1]), .C(raw_x_0), .D(n41438), .Z(bypass_data_0_31__N_872[1])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam bypass_data_0_31__I_15_i2_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 mux_683_i10_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[9]), .D(left_shift_result[9]), .Z(n1826[9])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i10_4_lut_4_lut.init = 16'hd1c0;
    PFUMX bypass_data_0_31__I_14_i16 (.BLUT(bypass_data_0_31__N_1002[15]), 
          .ALUT(bypass_data_0_31__N_872[15]), .C0(n39363), .Z(bypass_data_0[15])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_683_i2_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[1]), .D(left_shift_result[1]), .Z(n1826[1])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i2_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_683_i23_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[22]), .D(left_shift_result[22]), .Z(n1826[22])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i23_4_lut_4_lut.init = 16'hd1c0;
    FD1S3AX operand_w_i15 (.D(operand_w_31__N_840[15]), .CK(w_clk_cpu), 
            .Q(operand_w[15])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i15.GSR = "ENABLED";
    LUT4 mux_683_i18_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[17]), .D(left_shift_result[17]), .Z(n1826[17])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i18_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_683_i14_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[13]), .D(left_shift_result[13]), .Z(n1826[13])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i14_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_683_i7_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[6]), .D(left_shift_result[6]), .Z(n1826[6])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i7_4_lut_4_lut.init = 16'hd1c0;
    LUT4 valid_d_I_0_757_2_lut_rep_288_4_lut (.A(instruction_d[15]), .B(n42722), 
         .C(n41397), .D(valid_d), .Z(n41375)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(D))+!A (B+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1544[36:105])
    defparam valid_d_I_0_757_2_lut_rep_288_4_lut.init = 16'h3b00;
    FD1P3AX operand_m_i0_i4 (.D(x_result[4]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(operand_m[4])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i4.GSR = "ENABLED";
    LUT4 i38036_2_lut (.A(m_result_sel_compare_m), .B(m_result_sel_shift_m), 
         .Z(n39334)) /* synthesis lut_function=(A+!(B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1627[18] 1631[27])
    defparam i38036_2_lut.init = 16'hbbbb;
    FD1P3AX operand_m_i0_i3 (.D(x_result[3]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(operand_m[3])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i3.GSR = "ENABLED";
    LUT4 bypass_data_1_31__I_16_i13_3_lut (.A(m_result[12]), .B(x_result[12]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i13_3_lut.init = 16'hcaca;
    LUT4 mux_52_i13_3_lut (.A(reg_data_1[12]), .B(w_result[12]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i13_3_lut.init = 16'hcaca;
    LUT4 bypass_data_1_31__I_16_i12_3_lut (.A(m_result[11]), .B(x_result[11]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i12_3_lut.init = 16'hcaca;
    LUT4 mux_52_i12_3_lut (.A(reg_data_1[11]), .B(w_result[11]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i12_3_lut.init = 16'hcaca;
    FD1S3AX operand_w_i14 (.D(operand_w_31__N_840[14]), .CK(w_clk_cpu), 
            .Q(operand_w[14])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i14.GSR = "ENABLED";
    LUT4 mux_683_i4_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[3]), .D(left_shift_result[3]), .Z(n1826[3])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i4_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_683_i31_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[30]), .D(left_shift_result[30]), .Z(n1826[30])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i31_4_lut_4_lut.init = 16'hd1c0;
    FD1P3AX operand_m_i0_i2 (.D(x_result[2]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(operand_m[2])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i2.GSR = "ENABLED";
    LUT4 bypass_data_1_31__I_16_i11_3_lut (.A(m_result[10]), .B(x_result[10]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i11_3_lut.init = 16'hcaca;
    LUT4 mux_683_i29_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[28]), .D(left_shift_result[28]), .Z(n1826[28])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i29_4_lut_4_lut.init = 16'hd1c0;
    FD1P3AX operand_m_i0_i1 (.D(x_result[1]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(operand_m[1])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_m_i0_i1.GSR = "ENABLED";
    FD1S3AX operand_w_i13 (.D(operand_w_31__N_840[13]), .CK(w_clk_cpu), 
            .Q(operand_w[13])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i13.GSR = "ENABLED";
    LUT4 mux_52_i11_3_lut (.A(reg_data_1[10]), .B(w_result[10]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i11_3_lut.init = 16'hcaca;
    LUT4 bypass_data_1_31__I_16_i10_3_lut (.A(m_result[9]), .B(x_result[9]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i10_3_lut.init = 16'hcaca;
    LUT4 mux_52_i10_3_lut (.A(reg_data_1[9]), .B(w_result[9]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i10_3_lut.init = 16'hcaca;
    CCU2D operand_0_x_31__I_0_29 (.A0(operand_1_x[9]), .B0(muliplicand[9]), 
          .C0(operand_1_x[8]), .D0(muliplicand[8]), .A1(operand_1_x[7]), 
          .B1(muliplicand[7]), .C1(operand_1_x[6]), .D1(muliplicand[6]), 
          .CIN(n36491), .COUT(n36492));
    defparam operand_0_x_31__I_0_29.INIT0 = 16'h9009;
    defparam operand_0_x_31__I_0_29.INIT1 = 16'h9009;
    defparam operand_0_x_31__I_0_29.INJECT1_0 = "YES";
    defparam operand_0_x_31__I_0_29.INJECT1_1 = "YES";
    LUT4 branch_predict_m_bdd_3_lut (.A(branch_predict_m), .B(condition_met_m), 
         .C(branch_predict_taken_m), .Z(n41147)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A ((C)+!B))) */ ;
    defparam branch_predict_m_bdd_3_lut.init = 16'h2c2c;
    LUT4 i1_4_lut_rep_341 (.A(LM32I_CYC_O), .B(LM32D_CYC_O), .C(stall_wb_load), 
         .D(n52), .Z(n41428)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1924[21] 1957[39])
    defparam i1_4_lut_rep_341.init = 16'hfefa;
    LUT4 bypass_data_1_31__I_16_i9_3_lut (.A(m_result[8]), .B(x_result[8]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i9_3_lut.init = 16'hcaca;
    LUT4 mux_52_i9_3_lut (.A(reg_data_1[8]), .B(w_result[8]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i9_3_lut.init = 16'hcaca;
    LUT4 bypass_data_1_31__I_16_i8_3_lut (.A(m_result[7]), .B(x_result[7]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i8_3_lut.init = 16'hcaca;
    LUT4 mux_683_i28_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[27]), .D(left_shift_result[27]), .Z(n1826[27])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i28_4_lut_4_lut.init = 16'hd1c0;
    PFUMX bypass_data_0_31__I_14_i17 (.BLUT(bypass_data_0_31__N_1002[16]), 
          .ALUT(bypass_data_0_31__N_872[16]), .C0(n39363), .Z(bypass_data_0[16])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 stall_m_I_0_1_lut_rep_323_4_lut (.A(LM32I_CYC_O), .B(LM32D_CYC_O), 
         .C(stall_wb_load), .D(n52), .Z(w_clk_cpu_enable_985)) /* synthesis lut_function=(!(A+(B (C+(D))+!B (C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1924[21] 1957[39])
    defparam stall_m_I_0_1_lut_rep_323_4_lut.init = 16'h0105;
    LUT4 mux_683_i26_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[25]), .D(left_shift_result[25]), .Z(n1826[25])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i26_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_683_i24_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[23]), .D(left_shift_result[23]), .Z(n1826[23])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i24_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_683_i21_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[20]), .D(left_shift_result[20]), .Z(n1826[20])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i21_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_683_i20_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[19]), .D(left_shift_result[19]), .Z(n1826[19])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i20_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_683_i17_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[16]), .D(left_shift_result[16]), .Z(n1826[16])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i17_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_683_i15_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[14]), .D(left_shift_result[14]), .Z(n1826[14])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i15_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_683_i13_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[12]), .D(left_shift_result[12]), .Z(n1826[12])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i13_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_683_i9_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[8]), .D(left_shift_result[8]), .Z(n1826[8])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i9_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_52_i8_3_lut (.A(reg_data_1[7]), .B(w_result[7]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i8_3_lut.init = 16'hcaca;
    LUT4 mux_683_i8_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[7]), .D(left_shift_result[7]), .Z(n1826[7])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i8_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_683_i6_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[5]), .D(left_shift_result[5]), .Z(n1826[5])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i6_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_683_i5_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[4]), .D(left_shift_result[4]), .Z(n1826[4])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i5_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(eret_x), .B(n41391), .C(n25705), 
         .D(csr_write_enable_x), .Z(n4_adj_3898)) /* synthesis lut_function=(A (B)+!A !((C+!(D))+!B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1984[19:54])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h8c88;
    LUT4 ie_I_110_3_lut_4_lut (.A(eret_x), .B(n41391), .C(eie), .D(ie_N_2822), 
         .Z(ie_N_2821)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1984[19:54])
    defparam ie_I_110_3_lut_4_lut.init = 16'hf780;
    FD1S3AX operand_w_i12 (.D(operand_w_31__N_840[12]), .CK(w_clk_cpu), 
            .Q(operand_w[12])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i12.GSR = "ENABLED";
    LUT4 mux_683_i3_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[2]), .D(left_shift_result[2]), .Z(n1826[2])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i3_4_lut_4_lut.init = 16'hd1c0;
    FD1S3AX operand_w_i11 (.D(operand_w_31__N_840[11]), .CK(w_clk_cpu), 
            .Q(operand_w[11])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i11.GSR = "ENABLED";
    LUT4 mux_683_i32_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[31]), .D(left_shift_result[31]), .Z(n1826[31])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i32_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_683_i30_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[29]), .D(left_shift_result[29]), .Z(n1826[29])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i30_4_lut_4_lut.init = 16'hd1c0;
    LUT4 bypass_data_1_31__I_16_i7_3_lut (.A(m_result[6]), .B(x_result[6]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i7_3_lut.init = 16'hcaca;
    LUT4 mux_52_i7_3_lut (.A(reg_data_1[6]), .B(w_result[6]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i7_3_lut.init = 16'hcaca;
    LUT4 mux_683_i27_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[26]), .D(left_shift_result[26]), .Z(n1826[26])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i27_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_683_i25_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[24]), .D(left_shift_result[24]), .Z(n1826[24])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i25_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_683_i22_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[21]), .D(left_shift_result[21]), .Z(n1826[21])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i22_4_lut_4_lut.init = 16'hd1c0;
    LUT4 bypass_data_1_31__I_16_i6_3_lut (.A(m_result[5]), .B(x_result[5]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i6_3_lut.init = 16'hcaca;
    LUT4 i21279_3_lut (.A(valid_w), .B(debug_exception_w), .C(non_debug_exception_w), 
         .Z(jtag_reg_d_7__N_505)) /* synthesis lut_function=(A (B+(C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1184[30:76])
    defparam i21279_3_lut.init = 16'ha8a8;
    LUT4 mux_52_i6_3_lut (.A(reg_data_1[5]), .B(w_result[5]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i6_3_lut.init = 16'hcaca;
    LUT4 csr_x_2__bdd_4_lut_38169 (.A(eba[17]), .B(csr_x[1]), .C(csr_x[3]), 
         .D(csr_x[0]), .Z(n40565)) /* synthesis lut_function=(!(A ((C)+!B)+!A ((C+(D))+!B))) */ ;
    defparam csr_x_2__bdd_4_lut_38169.init = 16'h080c;
    LUT4 bypass_data_1_31__I_16_i5_3_lut (.A(m_result[4]), .B(x_result[4]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i5_3_lut.init = 16'hcaca;
    PFUMX bypass_data_0_31__I_14_i18 (.BLUT(bypass_data_0_31__N_1002[17]), 
          .ALUT(bypass_data_0_31__N_872[17]), .C0(n39363), .Z(bypass_data_0[17])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_52_i5_3_lut (.A(reg_data_1[4]), .B(w_result[4]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i5_3_lut.init = 16'hcaca;
    LUT4 mux_683_i19_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[18]), .D(left_shift_result[18]), .Z(n1826[18])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i19_4_lut_4_lut.init = 16'hd1c0;
    LUT4 bypass_data_1_31__I_16_i4_3_lut (.A(m_result[3]), .B(x_result[3]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i4_3_lut.init = 16'hcaca;
    LUT4 mux_683_i16_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[15]), .D(left_shift_result[15]), .Z(n1826[15])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i16_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_683_i12_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[11]), .D(left_shift_result[11]), .Z(n1826[11])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i12_4_lut_4_lut.init = 16'hd1c0;
    LUT4 mux_465_i11_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[12]), .C(eba[12]), 
         .Z(n41553)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i11_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    PFUMX i23_adj_371 (.BLUT(n3_adj_3815), .ALUT(n7_adj_3792), .C0(csr_x[3]), 
          .Z(n10_adj_3895));
    FD1S3AX operand_w_i10 (.D(operand_w_31__N_840[10]), .CK(w_clk_cpu), 
            .Q(operand_w[10])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i10.GSR = "ENABLED";
    LUT4 mux_683_i11_4_lut_4_lut (.A(m_result_sel_compare_m), .B(raw_x_1), 
         .C(n1253[10]), .D(left_shift_result[10]), .Z(n1826[10])) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam mux_683_i11_4_lut_4_lut.init = 16'hd1c0;
    FD1S3AX operand_w_i9 (.D(operand_w_31__N_840[9]), .CK(w_clk_cpu), .Q(operand_w[9])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i9.GSR = "ENABLED";
    FD1P3IX valid_d_618 (.D(valid_d_N_1264), .SP(w_clk_cpu_enable_638), 
            .CD(branch_taken_m), .CK(w_clk_cpu), .Q(valid_d));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2264[5] 2299[8])
    defparam valid_d_618.GSR = "ENABLED";
    LUT4 mux_52_i4_3_lut (.A(reg_data_1[3]), .B(w_result[3]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i4_3_lut.init = 16'hcaca;
    LUT4 bypass_data_1_31__I_16_i3_3_lut (.A(m_result[2]), .B(x_result[2]), 
         .C(raw_x_1), .Z(bypass_data_1_31__N_904[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1531[10] 1534[36])
    defparam bypass_data_1_31__I_16_i3_3_lut.init = 16'hcaca;
    PFUMX bypass_data_0_31__I_14_i19 (.BLUT(bypass_data_0_31__N_1002[18]), 
          .ALUT(bypass_data_0_31__N_872[18]), .C0(n39363), .Z(bypass_data_0[18])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i20117_2_lut_2_lut_3_lut (.A(n41526), .B(non_debug_exception_x_N_1357), 
         .C(n41428), .Z(n22503)) /* synthesis lut_function=(!(A (C)+!A ((C)+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam i20117_2_lut_2_lut_3_lut.init = 16'h0e0e;
    LUT4 mux_52_i3_3_lut (.A(reg_data_1[2]), .B(w_result[2]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i3_3_lut.init = 16'hcaca;
    PFUMX bypass_data_0_31__I_14_i20 (.BLUT(bypass_data_0_31__N_1002[19]), 
          .ALUT(bypass_data_0_31__N_872[19]), .C0(n39363), .Z(bypass_data_0[19])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 csr_x_2__bdd_4_lut_38547 (.A(deba[17]), .B(csr_x[1]), .C(csr_x[3]), 
         .D(csr_x[0]), .Z(n40566)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam csr_x_2__bdd_4_lut_38547.init = 16'h2000;
    LUT4 mux_465_i11_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[12]), .C(branch_target_x[12]), 
         .Z(n41552)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i11_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    FD1S3AX operand_w_i8 (.D(operand_w_31__N_840[8]), .CK(w_clk_cpu), .Q(operand_w[8])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i8.GSR = "ENABLED";
    LUT4 mux_52_i2_3_lut (.A(reg_data_1[1]), .B(w_result[1]), .C(raw_w_1), 
         .Z(bypass_data_1_31__N_1034[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1534[9:36])
    defparam mux_52_i2_3_lut.init = 16'hcaca;
    PFUMX bypass_data_0_31__I_14_i21 (.BLUT(bypass_data_0_31__N_1002[20]), 
          .ALUT(bypass_data_0_31__N_872[20]), .C0(n39363), .Z(bypass_data_0[20])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_2_lut_3_lut (.A(n41526), .B(non_debug_exception_x_N_1357), .C(write_idx_x[4]), 
         .Z(write_idx_m_4__N_1152[4])) /* synthesis lut_function=(A+(B+(C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    CCU2D operand_0_x_31__I_0_27 (.A0(operand_1_x[13]), .B0(muliplicand[13]), 
          .C0(operand_1_x[12]), .D0(muliplicand[12]), .A1(operand_1_x[11]), 
          .B1(muliplicand[11]), .C1(operand_1_x[10]), .D1(muliplicand[10]), 
          .CIN(n36490), .COUT(n36491));
    defparam operand_0_x_31__I_0_27.INIT0 = 16'h9009;
    defparam operand_0_x_31__I_0_27.INIT1 = 16'h9009;
    defparam operand_0_x_31__I_0_27.INJECT1_0 = "YES";
    defparam operand_0_x_31__I_0_27.INJECT1_1 = "YES";
    PFUMX i23_adj_372 (.BLUT(n3_adj_3814), .ALUT(n7_adj_3791), .C0(csr_x[3]), 
          .Z(n10_adj_3860));
    PFUMX bypass_data_0_31__I_14_i22 (.BLUT(bypass_data_0_31__N_1002[21]), 
          .ALUT(bypass_data_0_31__N_872[21]), .C0(n39363), .Z(bypass_data_0[21])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i1_2_lut_3_lut_adj_373 (.A(n41526), .B(non_debug_exception_x_N_1357), 
         .C(write_idx_x[2]), .Z(write_idx_m_4__N_1152[2])) /* synthesis lut_function=(A+(B+(C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam i1_2_lut_3_lut_adj_373.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_adj_374 (.A(n41526), .B(non_debug_exception_x_N_1357), 
         .C(write_idx_x[3]), .Z(write_idx_m_4__N_1152[3])) /* synthesis lut_function=(A+(B+(C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam i1_2_lut_3_lut_adj_374.init = 16'hfefe;
    PFUMX bypass_data_0_31__I_14_i23 (.BLUT(bypass_data_0_31__N_1002[22]), 
          .ALUT(bypass_data_0_31__N_872[22]), .C0(n39363), .Z(bypass_data_0[22])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX i23_adj_375 (.BLUT(n3_adj_3813), .ALUT(n7_adj_3790), .C0(csr_x[3]), 
          .Z(n10_adj_3881));
    FD1P3IX data_bus_error_exception_m_657 (.D(data_bus_error_exception), 
            .SP(w_clk_cpu_enable_711), .CD(n22524), .CK(w_clk_cpu), .Q(data_bus_error_exception_m));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam data_bus_error_exception_m_657.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_376 (.A(n41526), .B(non_debug_exception_x_N_1357), 
         .C(write_idx_x[1]), .Z(write_idx_m_4__N_1152[1])) /* synthesis lut_function=(A+(B+(C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam i1_2_lut_3_lut_adj_376.init = 16'hfefe;
    FD1S3AX operand_w_i7 (.D(operand_w_31__N_840[7]), .CK(w_clk_cpu), .Q(operand_w[7])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i7.GSR = "ENABLED";
    LUT4 i28961_2_lut_3_lut (.A(n41526), .B(non_debug_exception_x_N_1357), 
         .C(write_enable_x), .Z(write_enable_m_N_1313)) /* synthesis lut_function=(A+(B+(C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam i28961_2_lut_3_lut.init = 16'hfefe;
    LUT4 i2_4_lut_4_lut (.A(n25722), .B(n41387), .C(w_clk_cpu_enable_958), 
         .D(n25724), .Z(n38840)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1980[22:60])
    defparam i2_4_lut_4_lut.init = 16'h0080;
    FD1P3AX write_idx_m_i0_i4 (.D(write_idx_m_4__N_1152[4]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(write_idx_m[4])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_m_i0_i4.GSR = "ENABLED";
    PFUMX i23_adj_377 (.BLUT(n3_adj_3798), .ALUT(n7_adj_3789), .C0(csr_x[3]), 
          .Z(n10_adj_3891));
    LUT4 mux_465_i12_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[13]), .C(eba[13]), 
         .Z(n41556)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i12_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    FD1S3AX operand_w_i6 (.D(operand_w_31__N_840[6]), .CK(w_clk_cpu), .Q(operand_w[6])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i6.GSR = "ENABLED";
    FD1P3AX write_idx_m_i0_i3 (.D(write_idx_m_4__N_1152[3]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(write_idx_m[3])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_m_i0_i3.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_415 (.A(csr_x[3]), .B(csr_x[4]), .Z(n41502)) /* synthesis lut_function=((B)+!A) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2132[5:19])
    defparam i1_2_lut_rep_415.init = 16'hdddd;
    PFUMX bypass_data_0_31__I_14_i24 (.BLUT(bypass_data_0_31__N_1002[23]), 
          .ALUT(bypass_data_0_31__N_872[23]), .C0(n39363), .Z(bypass_data_0[23])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX bypass_data_0_31__I_14_i25 (.BLUT(bypass_data_0_31__N_1002[24]), 
          .ALUT(bypass_data_0_31__N_872[24]), .C0(n39363), .Z(bypass_data_0[24])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 i2_3_lut_rep_416 (.A(csr_x[2]), .B(csr_x[4]), .C(csr_x[1]), .Z(n41503)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i2_3_lut_rep_416.init = 16'h2020;
    LUT4 valid_f_I_0_2_lut_3_lut_4_lut (.A(valid_d), .B(n41394), .C(valid_f), 
         .D(branch_taken_m), .Z(valid_d_N_1264)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1690[20] 1692[7])
    defparam valid_f_I_0_2_lut_3_lut_4_lut.init = 16'h0070;
    FD1S3AX operand_w_i5 (.D(operand_w_31__N_840[5]), .CK(w_clk_cpu), .Q(operand_w[5])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i5.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_370_4_lut (.A(csr_x[2]), .B(csr_x[4]), .C(csr_x[1]), 
         .D(csr_x[3]), .Z(n41457)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i1_2_lut_rep_370_4_lut.init = 16'h0020;
    LUT4 i34124_2_lut_rep_417 (.A(pc_d[2]), .B(instruction_d[0]), .Z(n41504)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i34124_2_lut_rep_417.init = 16'h6666;
    LUT4 mux_389_i1_3_lut_4_lut (.A(pc_d[2]), .B(instruction_d[0]), .C(n22224), 
         .D(bypass_data_0[2]), .Z(branch_target_x_31__N_1122[0])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam mux_389_i1_3_lut_4_lut.init = 16'hf606;
    FD1P3AX write_idx_m_i0_i2 (.D(write_idx_m_4__N_1152[2]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(write_idx_m[2])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_m_i0_i2.GSR = "ENABLED";
    CCU2D operand_0_x_31__I_0_19 (.A0(operand_1_x[29]), .B0(muliplicand[29]), 
          .C0(operand_1_x[28]), .D0(muliplicand[28]), .A1(operand_1_x[27]), 
          .B1(muliplicand[27]), .C1(operand_1_x[26]), .D1(muliplicand[26]), 
          .CIN(n36486), .COUT(n36487));
    defparam operand_0_x_31__I_0_19.INIT0 = 16'h9009;
    defparam operand_0_x_31__I_0_19.INIT1 = 16'h9009;
    defparam operand_0_x_31__I_0_19.INJECT1_0 = "YES";
    defparam operand_0_x_31__I_0_19.INJECT1_1 = "YES";
    LUT4 i37805_2_lut (.A(write_idx_m[3]), .B(read_idx_1_d[3]), .Z(n39886)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(472[26:38])
    defparam i37805_2_lut.init = 16'h6666;
    FD1S3AX operand_w_i4 (.D(operand_w_31__N_840[4]), .CK(w_clk_cpu), .Q(operand_w[4])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i4.GSR = "ENABLED";
    LUT4 mux_465_i12_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[13]), .C(branch_target_x[13]), 
         .Z(n41555)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i12_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 i1_2_lut_rep_420 (.A(branch_predict_taken_m), .B(branch_predict_m), 
         .Z(n41507)) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1680[13] 1683[7])
    defparam i1_2_lut_rep_420.init = 16'h8888;
    LUT4 i2_4_lut_adj_378 (.A(write_idx_m[0]), .B(write_idx_m[2]), .C(read_idx_1_d[0]), 
         .D(read_idx_1_d[2]), .Z(n6)) /* synthesis lut_function=(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(472[26:38])
    defparam i2_4_lut_adj_378.init = 16'h8421;
    FD1P3AX write_idx_m_i0_i1 (.D(write_idx_m_4__N_1152[1]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(write_idx_m[1])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_m_i0_i1.GSR = "ENABLED";
    FD1P3AX m_result_sel_shift_x_632 (.D(m_result_sel_shift_d), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(m_result_sel_shift_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam m_result_sel_shift_x_632.GSR = "ENABLED";
    FD1P3AX w_result_sel_mul_x_634 (.D(w_result_sel_mul_d), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(w_result_sel_mul_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam w_result_sel_mul_x_634.GSR = "ENABLED";
    FD1P3AX x_bypass_enable_x_635 (.D(x_bypass_enable_d), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(x_bypass_enable_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam x_bypass_enable_x_635.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_372_3_lut (.A(branch_predict_taken_m), .B(branch_predict_m), 
         .C(condition_met_m), .Z(n41459)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1680[13] 1683[7])
    defparam i1_2_lut_rep_372_3_lut.init = 16'h0808;
    FD1P3AX m_bypass_enable_x_636 (.D(m_bypass_enable_d), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(m_bypass_enable_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam m_bypass_enable_x_636.GSR = "ENABLED";
    FD1S3AX operand_w_i3 (.D(operand_w_31__N_840[3]), .CK(w_clk_cpu), .Q(operand_w[3])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i3.GSR = "ENABLED";
    LUT4 mux_19150_i8_3_lut_4_lut (.A(size_x[1]), .B(condition_x[0]), .C(muliplicand[7]), 
         .D(muliplicand[15]), .Z(n21411[21])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_19150_i8_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_19150_i7_3_lut_4_lut (.A(size_x[1]), .B(condition_x[0]), .C(muliplicand[7]), 
         .D(muliplicand[14]), .Z(n21411[6])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_19150_i7_3_lut_4_lut.init = 16'hfe10;
    LUT4 i37222_3_lut_4_lut (.A(cmp_zero), .B(condition_x[0]), .C(size_x[1]), 
         .D(adder_carry_n_x), .Z(n39776)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !(C+(D)))) */ ;
    defparam i37222_3_lut_4_lut.init = 16'h7770;
    LUT4 mux_19150_i6_3_lut_4_lut (.A(size_x[1]), .B(condition_x[0]), .C(muliplicand[7]), 
         .D(muliplicand[13]), .Z(n21411[5])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_19150_i6_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_19150_i5_3_lut_4_lut (.A(size_x[1]), .B(condition_x[0]), .C(muliplicand[7]), 
         .D(muliplicand[12]), .Z(n21411[4])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_19150_i5_3_lut_4_lut.init = 16'hfe10;
    FD1P3AX write_enable_x_637 (.D(write_enable_N_1809), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(write_enable_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_enable_x_637.GSR = "ENABLED";
    FD1P3AX size_x_i0_i1 (.D(size_d[1]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(size_x[1])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam size_x_i0_i1.GSR = "ENABLED";
    FD1S3AX operand_w_i2 (.D(operand_w_31__N_840[2]), .CK(w_clk_cpu), .Q(operand_w[2])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i2.GSR = "ENABLED";
    LUT4 mux_19150_i4_3_lut_4_lut (.A(size_x[1]), .B(condition_x[0]), .C(muliplicand[7]), 
         .D(muliplicand[11]), .Z(n21411[3])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_19150_i4_3_lut_4_lut.init = 16'hfe10;
    LUT4 i37809_2_lut (.A(write_idx_m[4]), .B(read_idx_1_d[4]), .Z(n39890)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(472[26:38])
    defparam i37809_2_lut.init = 16'h6666;
    FD1P3AX adder_op_x_n_645 (.D(adder_op_d_N_1339), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(adder_op_x_n));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam adder_op_x_n_645.GSR = "ENABLED";
    CCU2D operand_0_x_31__I_0_25 (.A0(operand_1_x[17]), .B0(muliplicand[17]), 
          .C0(operand_1_x[16]), .D0(muliplicand[16]), .A1(operand_1_x[15]), 
          .B1(muliplicand[15]), .C1(operand_1_x[14]), .D1(muliplicand[14]), 
          .CIN(n36489), .COUT(n36490));
    defparam operand_0_x_31__I_0_25.INIT0 = 16'h9009;
    defparam operand_0_x_31__I_0_25.INIT1 = 16'h9009;
    defparam operand_0_x_31__I_0_25.INJECT1_0 = "YES";
    defparam operand_0_x_31__I_0_25.INJECT1_1 = "YES";
    LUT4 mux_19150_i3_3_lut_4_lut (.A(size_x[1]), .B(condition_x[0]), .C(muliplicand[7]), 
         .D(muliplicand[10]), .Z(n21411[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_19150_i3_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_19150_i2_3_lut_4_lut (.A(size_x[1]), .B(condition_x[0]), .C(muliplicand[7]), 
         .D(muliplicand[9]), .Z(n21411[1])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_19150_i2_3_lut_4_lut.init = 16'hfe10;
    LUT4 mux_19150_i1_3_lut_4_lut (.A(size_x[1]), .B(condition_x[0]), .C(muliplicand[7]), 
         .D(muliplicand[8]), .Z(n21411[0])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;
    defparam mux_19150_i1_3_lut_4_lut.init = 16'hfe10;
    FD1P3AX branch_predict_x_649 (.D(branch_predict_d), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_predict_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_predict_x_649.GSR = "ENABLED";
    FD1P3AX branch_predict_taken_x_650 (.D(n41394), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(branch_predict_taken_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_predict_taken_x_650.GSR = "ENABLED";
    FD1S3IX operand_w_i1 (.D(n41438), .CK(w_clk_cpu), .CD(n24298), .Q(operand_w[1])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam operand_w_i1.GSR = "ENABLED";
    FD1P3AX eba_i8_i31 (.D(operand_1_x[31]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[31])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i31.GSR = "ENABLED";
    FD1P3IX branch_target_m_i2_i2 (.D(branch_target_x[2]), .SP(w_clk_cpu_enable_972), 
            .CD(n22503), .CK(w_clk_cpu), .Q(branch_target_m[2])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i2.GSR = "ENABLED";
    LUT4 i2_1_lut (.A(cycles_5__N_2495), .Z(mc_stall_request_x)) /* synthesis lut_function=(!(A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2285[14] 2286[34])
    defparam i2_1_lut.init = 16'h5555;
    LUT4 i2_4_lut_adj_379 (.A(divide_by_zero_x), .B(valid_x), .C(n23893), 
         .D(n31661), .Z(non_debug_exception_x_N_1357)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(377[5:12])
    defparam i2_4_lut_adj_379.init = 16'hfefa;
    FD1P3IX valid_x_619 (.D(n41387), .SP(w_clk_cpu_enable_697), .CD(n26126), 
            .CK(w_clk_cpu), .Q(valid_x)) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2264[5] 2299[8])
    defparam valid_x_619.GSR = "ENABLED";
    PFUMX x_result_31__I_0_i4 (.BLUT(x_result_31__N_1066[3]), .ALUT(x_result_31__N_616[3]), 
          .C0(n39459), .Z(x_result[3])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_389_i7_3_lut (.A(branch_target_d[8]), .B(bypass_data_0[8]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i7_3_lut.init = 16'hcaca;
    LUT4 mux_389_i6_3_lut (.A(branch_target_d[7]), .B(bypass_data_0[7]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i6_3_lut.init = 16'hcaca;
    LUT4 m_result_31__I_0_i17_3_lut (.A(m_result[16]), .B(operand_w_31__N_1187[16]), 
         .C(n42746), .Z(operand_w_31__N_840[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i17_3_lut.init = 16'hcaca;
    PFUMX x_result_31__I_0_i9 (.BLUT(sext_result_x[8]), .ALUT(x_result_31__N_616[8]), 
          .C0(n39497), .Z(x_result[8])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX eret_x_654 (.D(eret_d), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(eret_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam eret_x_654.GSR = "ENABLED";
    FD1P3AX bret_x_655 (.D(bret_d), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(bret_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam bret_x_655.GSR = "ENABLED";
    FD1P3AX bus_error_x_656 (.D(bus_error_d), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(bus_error_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam bus_error_x_656.GSR = "ENABLED";
    FD1P3AX csr_write_enable_x_658 (.D(n41406), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(csr_write_enable_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam csr_write_enable_x_658.GSR = "ENABLED";
    LUT4 write_idx_x_1__bdd_4_lut (.A(write_idx_x[1]), .B(read_idx_0_d[1]), 
         .C(read_idx_0_d[3]), .D(write_idx_x[3]), .Z(n40464)) /* synthesis lut_function=(A (B (C (D)+!C !(D)))+!A !(B+!(C (D)+!C !(D)))) */ ;
    defparam write_idx_x_1__bdd_4_lut.init = 16'h9009;
    FD1P3AX store_x_641 (.D(store_d), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(store_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_x_641.GSR = "ENABLED";
    FD1P3AX eba_i8_i30 (.D(operand_1_x[30]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[30])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i30.GSR = "ENABLED";
    LUT4 i1_3_lut_rep_345 (.A(csr_x[0]), .B(csr_x[3]), .C(n41503), .Z(n41432)) /* synthesis lut_function=(A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i1_3_lut_rep_345.init = 16'h8080;
    LUT4 i1_2_lut_adj_380 (.A(bus_error_x), .B(scall_x), .Z(n31661)) /* synthesis lut_function=(A+(B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(377[5:12])
    defparam i1_2_lut_adj_380.init = 16'heeee;
    LUT4 i1_2_lut_4_lut_adj_381 (.A(csr_x[0]), .B(csr_x[3]), .C(n41503), 
         .D(jrx_csr_read_data[3]), .Z(n36690)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i1_2_lut_4_lut_adj_381.init = 16'h8000;
    LUT4 mux_389_i5_3_lut (.A(branch_target_d[6]), .B(bypass_data_0[6]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i5_3_lut.init = 16'hcaca;
    LUT4 mux_389_i4_3_lut (.A(branch_target_d[5]), .B(bypass_data_0[5]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i4_3_lut.init = 16'hcaca;
    LUT4 mux_389_i3_3_lut (.A(branch_target_d[4]), .B(bypass_data_0[4]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i3_3_lut.init = 16'hcaca;
    PFUMX x_result_31__I_0_i10 (.BLUT(sext_result_x[9]), .ALUT(x_result_31__N_616[9]), 
          .C0(n39497), .Z(x_result[9])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_389_i2_3_lut (.A(branch_target_d[3]), .B(bypass_data_0[3]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i2_3_lut.init = 16'hcaca;
    LUT4 i21282_2_lut (.A(data_bus_error_exception), .B(reset_exception), 
         .Z(n23893)) /* synthesis lut_function=(A+(B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1829[10] 1864[33])
    defparam i21282_2_lut.init = 16'heeee;
    PFUMX x_result_31__I_0_i11 (.BLUT(sext_result_x[10]), .ALUT(x_result_31__N_616[10]), 
          .C0(n39497), .Z(x_result[10])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX m_bypass_enable_m_665 (.D(m_bypass_enable_x), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(m_bypass_enable_m));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam m_bypass_enable_m_665.GSR = "ENABLED";
    PFUMX i23_adj_382 (.BLUT(n3_adj_3812), .ALUT(n7_adj_3779), .C0(csr_x[3]), 
          .Z(n10_adj_3845));
    FD1P3IX w_result_sel_mul_m_664 (.D(w_result_sel_mul_x), .SP(w_clk_cpu_enable_711), 
            .CD(n22503), .CK(w_clk_cpu), .Q(w_result_sel_mul_m));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam w_result_sel_mul_m_664.GSR = "ENABLED";
    FD1P3AX adder_op_x_644 (.D(n41376), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(adder_op_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam adder_op_x_644.GSR = "ENABLED";
    FD1P3AX branch_m_666 (.D(branch_x), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(branch_m));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_m_666.GSR = "ENABLED";
    FD1P3AX branch_predict_m_667 (.D(branch_predict_x), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(branch_predict_m));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_predict_m_667.GSR = "ENABLED";
    FD1P3AX branch_predict_taken_m_668 (.D(branch_predict_taken_x), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(branch_predict_taken_m));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_predict_taken_m_668.GSR = "ENABLED";
    FD1P3AX eba_i8_i29 (.D(operand_1_x[29]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[29])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i29.GSR = "ENABLED";
    LUT4 mux_75_i27_3_lut (.A(logic_result_x[26]), .B(mc_result_x[26]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i27_3_lut.init = 16'hcaca;
    LUT4 mux_465_i7_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[8]), .C(eba[8]), 
         .Z(n41541)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i7_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 i1_2_lut_rep_425 (.A(valid_m), .B(n42746), .Z(n41512)) /* synthesis lut_function=(!((B)+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(746[5:16])
    defparam i1_2_lut_rep_425.init = 16'h2222;
    LUT4 i1_2_lut_rep_285_3_lut_3_lut_4_lut (.A(valid_m), .B(n42746), .C(store_m), 
         .D(n41428), .Z(n41372)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(746[5:16])
    defparam i1_2_lut_rep_285_3_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(valid_m), .B(n42746), .C(n41493), 
         .D(LM32D_CYC_O), .Z(n4_adj_3899)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(746[5:16])
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_rep_426 (.A(load_m), .B(store_m), .Z(n41513)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_426.init = 16'heeee;
    PFUMX x_result_31__I_0_i12 (.BLUT(sext_result_x[11]), .ALUT(x_result_31__N_616[11]), 
          .C0(n39497), .Z(x_result[11])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX load_m_670 (.D(load_x), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(load_m));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam load_m_670.GSR = "ENABLED";
    LUT4 mux_465_i13_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[14]), .C(eba[14]), 
         .Z(n41562)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i13_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    PFUMX x_result_31__I_0_i13 (.BLUT(sext_result_x[12]), .ALUT(x_result_31__N_616[12]), 
          .C0(n39497), .Z(x_result[12])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 operand_m_31__I_0_704_i2_3_lut_rep_351 (.A(operand_m[1]), .B(shifter_result_m[1]), 
         .C(m_result_sel_shift_m), .Z(n41438)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1629[18] 1631[27])
    defparam operand_m_31__I_0_704_i2_3_lut_rep_351.init = 16'hcaca;
    PFUMX x_result_31__I_0_i14 (.BLUT(sext_result_x[13]), .ALUT(x_result_31__N_616[13]), 
          .C0(n39497), .Z(x_result[13])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX store_m_671 (.D(store_x), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(store_m));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam store_m_671.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_383 (.A(load_m), .B(store_m), .C(load_x), 
         .Z(n52)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_3_lut_adj_383.init = 16'hfefe;
    FD1P3AX eba_i8_i28 (.D(operand_1_x[28]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[28])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i28.GSR = "ENABLED";
    FD1P3AX eba_i8_i27 (.D(operand_1_x[27]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[27])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i27.GSR = "ENABLED";
    PFUMX x_result_31__I_0_i15 (.BLUT(sext_result_x[14]), .ALUT(x_result_31__N_616[14]), 
          .C0(n39497), .Z(x_result[14])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 operand_w_31__I_0_i32_3_lut (.A(operand_w[31]), .B(multiplier_result_w[31]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i32_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_384 (.A(n41531), .B(n39086), .C(n3_adj_3806), .D(n39126), 
         .Z(raw_w_1)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_384.init = 16'h0002;
    LUT4 operand_w_31__I_0_i31_3_lut (.A(operand_w[30]), .B(multiplier_result_w[30]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i31_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i18_3_lut (.A(operand_w[17]), .B(multiplier_result_w[17]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i18_3_lut.init = 16'hcaca;
    LUT4 mux_465_i13_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[14]), .C(branch_target_x[14]), 
         .Z(n41561)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i13_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    PFUMX x_result_31__I_0_i1 (.BLUT(x_result_31__N_1066[0]), .ALUT(x_result_31__N_616[0]), 
          .C0(n39459), .Z(x_result[0])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 operand_w_31__I_0_i17_3_lut (.A(operand_w[16]), .B(multiplier_result_w[16]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i17_3_lut.init = 16'hcaca;
    FD1P3AX eba_i8_i26 (.D(operand_1_x[26]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[26])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i26.GSR = "ENABLED";
    LUT4 mux_465_i15_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[16]), .C(eba[16]), 
         .Z(n41568)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i15_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    FD1P3AX eba_i8_i25 (.D(operand_1_x[25]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[25])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i25.GSR = "ENABLED";
    PFUMX x_result_31__I_0_i5 (.BLUT(x_result_31__N_1066[4]), .ALUT(x_result_31__N_616[4]), 
          .C0(n39459), .Z(x_result[4])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_19174_i15_3_lut (.A(pc_m[16]), .B(memop_pc_w[16]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i15_3_lut.init = 16'hcaca;
    PFUMX x_result_31__I_0_i6 (.BLUT(x_result_31__N_1066[5]), .ALUT(x_result_31__N_616[5]), 
          .C0(n39459), .Z(x_result[5])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX eba_i8_i24 (.D(operand_1_x[24]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[24])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i24.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_385 (.A(valid_m), .B(write_enable_m), .Z(n34433)) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2264[5] 2299[8])
    defparam i1_2_lut_adj_385.init = 16'h8888;
    PFUMX x_result_31__I_0_i7 (.BLUT(x_result_31__N_1066[6]), .ALUT(x_result_31__N_616[6]), 
          .C0(n39459), .Z(x_result[6])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX eba_i8_i23 (.D(operand_1_x[23]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[23])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i23.GSR = "ENABLED";
    LUT4 mux_389_i30_3_lut (.A(branch_target_d[31]), .B(bypass_data_0[31]), 
         .C(n22224), .Z(branch_target_x_31__N_1122[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2429[35:104])
    defparam mux_389_i30_3_lut.init = 16'hcaca;
    PFUMX x_result_31__I_0_i8 (.BLUT(x_result_31__N_1066[7]), .ALUT(x_result_31__N_616[7]), 
          .C0(n39459), .Z(x_result[7])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX i38573 (.BLUT(n41543), .ALUT(n41544), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[7]));
    LUT4 mux_20532_i5_3_lut (.A(n23056), .B(n23088), .C(read_idx_0_d[4]), 
         .Z(n23116[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i5_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i16_3_lut (.A(operand_w[15]), .B(multiplier_result_w[15]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i16_3_lut.init = 16'hcaca;
    PFUMX x_result_31__I_0_i16 (.BLUT(x_result_31__N_1066[15]), .ALUT(x_result_31__N_616[15]), 
          .C0(n39459), .Z(x_result[15])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX eba_i8_i22 (.D(operand_1_x[22]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[22])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i22.GSR = "ENABLED";
    LUT4 mux_465_i15_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[16]), .C(branch_target_x[16]), 
         .Z(n41567)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i15_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    FD1P3AX eba_i8_i21 (.D(operand_1_x[21]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[21])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i21.GSR = "ENABLED";
    PFUMX x_result_31__I_0_i17 (.BLUT(x_result_31__N_1066[16]), .ALUT(x_result_31__N_616[16]), 
          .C0(n39459), .Z(x_result[16])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_20532_i6_3_lut (.A(n23057), .B(n23089), .C(read_idx_0_d[4]), 
         .Z(n23116[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i6_3_lut.init = 16'hcaca;
    PFUMX x_result_31__I_0_i18 (.BLUT(x_result_31__N_1066[17]), .ALUT(x_result_31__N_616[17]), 
          .C0(n39459), .Z(x_result[17])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX i38571 (.BLUT(n41540), .ALUT(n41541), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[6]));
    LUT4 operand_w_31__I_0_i15_3_lut (.A(operand_w[14]), .B(multiplier_result_w[14]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i15_3_lut.init = 16'hcaca;
    FD1P3AX eba_i8_i20 (.D(operand_1_x[20]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[20])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i20.GSR = "ENABLED";
    FD1P3AX write_enable_m_672 (.D(write_enable_m_N_1313), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(write_enable_m));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_enable_m_672.GSR = "ENABLED";
    LUT4 operand_w_31__I_0_i14_3_lut (.A(operand_w[13]), .B(multiplier_result_w[13]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i14_3_lut.init = 16'hcaca;
    PFUMX x_result_31__I_0_i19 (.BLUT(x_result_31__N_1066[18]), .ALUT(x_result_31__N_616[18]), 
          .C0(n39459), .Z(x_result[18])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3IX exception_m_669_rep_465 (.D(exception_m_N_1355), .SP(w_clk_cpu_enable_972), 
            .CD(n31636), .CK(w_clk_cpu), .Q(n42746));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam exception_m_669_rep_465.GSR = "ENABLED";
    FD1P3AX eba_i8_i19 (.D(operand_1_x[19]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[19])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i19.GSR = "ENABLED";
    LUT4 mux_465_i16_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[17]), .C(eba[17]), 
         .Z(n41571)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i16_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    PFUMX x_result_31__I_0_i20 (.BLUT(x_result_31__N_1066[19]), .ALUT(x_result_31__N_616[19]), 
          .C0(n39459), .Z(x_result[19])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX eba_i8_i18 (.D(operand_1_x[18]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[18])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i18.GSR = "ENABLED";
    LUT4 i1_3_lut_adj_386 (.A(n41526), .B(non_debug_exception_x_N_1357), 
         .C(write_idx_x[0]), .Z(write_idx_m_4__N_1152[0])) /* synthesis lut_function=(!(A (B)+!A (B+!(C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(771[6:26])
    defparam i1_3_lut_adj_386.init = 16'h3232;
    FD1P3AX non_debug_exception_m_676 (.D(non_debug_exception_x_N_1357), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(non_debug_exception_m));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam non_debug_exception_m_676.GSR = "ENABLED";
    PFUMX x_result_31__I_0_i21 (.BLUT(x_result_31__N_1066[20]), .ALUT(x_result_31__N_616[20]), 
          .C0(n39459), .Z(x_result[20])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 operand_w_31__I_0_i13_3_lut (.A(operand_w[12]), .B(multiplier_result_w[12]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i13_3_lut.init = 16'hcaca;
    LUT4 mux_465_i16_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[17]), .C(branch_target_x[17]), 
         .Z(n41570)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i16_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    FD1P3AX eba_i8_i17 (.D(operand_1_x[17]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[17])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i17.GSR = "ENABLED";
    FD1P3AX eba_i8_i16 (.D(operand_1_x[16]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[16])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i16.GSR = "ENABLED";
    PFUMX x_result_31__I_0_i22 (.BLUT(x_result_31__N_1066[21]), .ALUT(x_result_31__N_616[21]), 
          .C0(n39459), .Z(x_result[21])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_465_i30_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[31]), .C(eba[31]), 
         .Z(n41574)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i30_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    PFUMX x_result_31__I_0_i23 (.BLUT(x_result_31__N_1066[22]), .ALUT(x_result_31__N_616[22]), 
          .C0(n39459), .Z(x_result[22])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX eba_i8_i15 (.D(operand_1_x[15]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[15])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i15.GSR = "ENABLED";
    LUT4 operand_w_31__I_0_i12_3_lut (.A(operand_w[11]), .B(multiplier_result_w[11]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 mux_465_i30_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[31]), .C(branch_target_x[31]), 
         .Z(n41573)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i30_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    PFUMX x_result_31__I_0_i24 (.BLUT(x_result_31__N_1066[23]), .ALUT(x_result_31__N_616[23]), 
          .C0(n39459), .Z(x_result[23])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX eba_i8_i14 (.D(operand_1_x[14]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[14])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i14.GSR = "ENABLED";
    PFUMX x_result_31__I_0_i25 (.BLUT(x_result_31__N_1066[24]), .ALUT(x_result_31__N_616[24]), 
          .C0(n39459), .Z(x_result[24])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX eba_i8_i13 (.D(operand_1_x[13]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[13])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i13.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut_3_lut (.A(n41474), .B(csr_x[1]), .C(csr_x[0]), 
         .Z(n38878)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_3_lut_4_lut_3_lut.init = 16'h1010;
    FD1P3AX eba_i8_i12 (.D(operand_1_x[12]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[12])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i12.GSR = "ENABLED";
    FD1S3AX write_idx_w_i0_rep_457 (.D(write_idx_m[0]), .CK(w_clk_cpu), 
            .Q(n42738)) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_w_i0_rep_457.GSR = "ENABLED";
    PFUMX x_result_31__I_0_i26 (.BLUT(x_result_31__N_1066[25]), .ALUT(x_result_31__N_616[25]), 
          .C0(n39459), .Z(x_result[25])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i27 (.BLUT(x_result_31__N_1066[26]), .ALUT(x_result_31__N_616[26]), 
          .C0(n39459), .Z(x_result[26])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1P3AX eba_i8_i11 (.D(operand_1_x[11]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[11])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i11.GSR = "ENABLED";
    FD1P3AX eba_i8_i10 (.D(operand_1_x[10]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[10])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i10.GSR = "ENABLED";
    LUT4 csr_x_2__bdd_4_lut_38548 (.A(eba[27]), .B(csr_x[1]), .C(csr_x[3]), 
         .D(csr_x[0]), .Z(n41319)) /* synthesis lut_function=(!(A ((C)+!B)+!A ((C+(D))+!B))) */ ;
    defparam csr_x_2__bdd_4_lut_38548.init = 16'h080c;
    FD1P3AX eba_i8_i9 (.D(operand_1_x[9]), .SP(eba_31__N_1101), .CK(w_clk_cpu), 
            .Q(eba[9])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2154[5] 2161[8])
    defparam eba_i8_i9.GSR = "ENABLED";
    FD1P3AX m_result_sel_shift_m_662_rep_455 (.D(m_result_sel_shift_x), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(n42736));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam m_result_sel_shift_m_662_rep_455.GSR = "ENABLED";
    PFUMX x_result_31__I_0_i28 (.BLUT(x_result_31__N_1066[27]), .ALUT(x_result_31__N_616[27]), 
          .C0(n39459), .Z(x_result[27])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    PFUMX x_result_31__I_0_i29 (.BLUT(x_result_31__N_1066[28]), .ALUT(x_result_31__N_616[28]), 
          .C0(n39459), .Z(x_result[28])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    FD1S3AX write_idx_w_i3_rep_453 (.D(write_idx_m[3]), .CK(w_clk_cpu), 
            .Q(n42734)) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_w_i3_rep_453.GSR = "ENABLED";
    PFUMX x_result_31__I_0_i30 (.BLUT(x_result_31__N_1066[29]), .ALUT(x_result_31__N_616[29]), 
          .C0(n39459), .Z(x_result[29])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 m_result_31__I_0_i20_3_lut (.A(m_result[19]), .B(operand_w_31__N_1187[19]), 
         .C(n42746), .Z(operand_w_31__N_840[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i20_3_lut.init = 16'hcaca;
    LUT4 csr_x_2__bdd_4_lut (.A(deba[27]), .B(csr_x[1]), .C(csr_x[3]), 
         .D(csr_x[0]), .Z(n41320)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam csr_x_2__bdd_4_lut.init = 16'h2000;
    FD1P3AX branch_target_m_i2_i31 (.D(branch_target_m_31__N_1157[29]), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(branch_target_m[31])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i31.GSR = "ENABLED";
    PFUMX x_result_31__I_0_i31 (.BLUT(x_result_31__N_1066[30]), .ALUT(x_result_31__N_616[30]), 
          .C0(n39459), .Z(x_result[30])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 mux_19174_i18_3_lut (.A(pc_m[19]), .B(memop_pc_w[19]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i18_3_lut.init = 16'hcaca;
    FD1S3AX write_idx_w_i2_rep_451 (.D(write_idx_m[2]), .CK(w_clk_cpu), 
            .Q(n42732)) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam write_idx_w_i2_rep_451.GSR = "ENABLED";
    PFUMX x_result_31__I_0_i32 (.BLUT(x_result_31__N_1066[31]), .ALUT(x_result_31__N_616[31]), 
          .C0(n39459), .Z(x_result[31])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    LUT4 operand_w_31__I_0_i2_3_lut (.A(operand_w[1]), .B(multiplier_result_w[1]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i2_3_lut.init = 16'hcaca;
    FD1P3AX branch_target_m_i2_i30 (.D(branch_target_m_31__N_1157[28]), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(branch_target_m[30])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i30.GSR = "ENABLED";
    FD1P3AX branch_target_m_i2_i29 (.D(branch_target_m_31__N_1157[27]), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(branch_target_m[29])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i29.GSR = "ENABLED";
    FD1P3AX branch_target_m_i2_i28 (.D(branch_target_m_31__N_1157[26]), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(branch_target_m[28])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i28.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_387 (.A(n9_adj_3900), .B(muliplicand[31]), .C(adder_result_x[31]), 
         .D(operand_1_x[31]), .Z(n24748)) /* synthesis lut_function=(!((B (C+!(D))+!B !((D)+!C))+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(713[6:14])
    defparam i1_4_lut_adj_387.init = 16'h2a02;
    LUT4 i1_2_lut_adj_388 (.A(cmp_zero), .B(condition_x[0]), .Z(n9_adj_3900)) /* synthesis lut_function=((B)+!A) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(713[6:14])
    defparam i1_2_lut_adj_388.init = 16'hdddd;
    LUT4 mux_465_i19_3_lut_4_lut_then_3_lut (.A(dc_re), .B(deba[20]), .C(eba[20]), 
         .Z(n41577)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i19_3_lut_4_lut_then_3_lut.init = 16'hd8d8;
    LUT4 mux_465_i19_3_lut_4_lut_else_3_lut (.A(n41526), .B(deba[20]), .C(branch_target_x[20]), 
         .Z(n41576)) /* synthesis lut_function=(A (B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1734[34] 1740[55])
    defparam mux_465_i19_3_lut_4_lut_else_3_lut.init = 16'hd8d8;
    LUT4 i20440_3_lut_4_lut (.A(n41531), .B(\counter[2] ), .C(n22999), 
         .D(write_idx_w[4]), .Z(n22877)) /* synthesis lut_function=(A (B ((D)+!C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2700[10] 2703[12])
    defparam i20440_3_lut_4_lut.init = 16'h8808;
    LUT4 i20437_3_lut_4_lut (.A(n41531), .B(\counter[2] ), .C(n22999), 
         .D(write_idx_w[4]), .Z(n22874)) /* synthesis lut_function=(!(((C (D))+!B)+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2700[10] 2703[12])
    defparam i20437_3_lut_4_lut.init = 16'h0888;
    FD1P3AX branch_target_m_i2_i27 (.D(branch_target_m_31__N_1157[25]), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(branch_target_m[27])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i27.GSR = "ENABLED";
    LUT4 mux_20532_i2_3_lut (.A(n23053), .B(n23085), .C(read_idx_0_d[4]), 
         .Z(n23116[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_389 (.A(n41531), .B(n39150), .C(n3_adj_3901), .D(n39082), 
         .Z(raw_w_0)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_389.init = 16'h0002;
    LUT4 i36603_4_lut (.A(write_idx_w[3]), .B(n42738), .C(read_idx_0_d[3]), 
         .D(read_idx_0_d[0]), .Z(n39150)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i36603_4_lut.init = 16'h7bde;
    LUT4 write_idx_w_4__I_0_748_i3_2_lut (.A(n42732), .B(read_idx_0_d[2]), 
         .Z(n3_adj_3901)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1487[18:47])
    defparam write_idx_w_4__I_0_748_i3_2_lut.init = 16'h6666;
    LUT4 i36536_4_lut (.A(write_idx_w[1]), .B(write_idx_w[4]), .C(read_idx_0_d[1]), 
         .D(read_idx_0_d[4]), .Z(n39082)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i36536_4_lut.init = 16'h7bde;
    LUT4 operand_w_31__I_0_i11_3_lut (.A(operand_w[10]), .B(multiplier_result_w[10]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 i3_4_lut_adj_390 (.A(valid_x), .B(n41408), .C(write_enable_x), 
         .D(n38827), .Z(raw_x_0)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2264[5] 2299[8])
    defparam i3_4_lut_adj_390.init = 16'h2000;
    LUT4 i2_4_lut_adj_391 (.A(write_idx_x[2]), .B(n4_adj_3902), .C(n40464), 
         .D(read_idx_0_d[2]), .Z(n38827)) /* synthesis lut_function=(A (B (C (D)))+!A !(((D)+!C)+!B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2264[5] 2299[8])
    defparam i2_4_lut_adj_391.init = 16'h8040;
    LUT4 i1_4_lut_adj_392 (.A(write_idx_x[0]), .B(write_idx_x[4]), .C(read_idx_0_d[0]), 
         .D(read_idx_0_d[4]), .Z(n4_adj_3902)) /* synthesis lut_function=(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2264[5] 2299[8])
    defparam i1_4_lut_adj_392.init = 16'h8421;
    LUT4 i37995_2_lut (.A(raw_x_0), .B(raw_m_0), .Z(n39363)) /* synthesis lut_function=(A+(B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1516[10] 1521[36])
    defparam i37995_2_lut.init = 16'heeee;
    FD1P3AX branch_target_m_i2_i26 (.D(branch_target_m_31__N_1157[24]), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(branch_target_m[26])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i26.GSR = "ENABLED";
    LUT4 debug_exception_w_I_0_2_lut_rep_385 (.A(debug_exception_w), .B(valid_w), 
         .Z(n41472)) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2007[30:82])
    defparam debug_exception_w_I_0_2_lut_rep_385.init = 16'h8888;
    LUT4 bie_I_115_3_lut_4_lut (.A(debug_exception_w), .B(valid_w), .C(ie), 
         .D(operand_1_x[2]), .Z(bie_N_2835)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2007[30:82])
    defparam bie_I_115_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_264_3_lut (.A(debug_exception_w), .B(valid_w), .C(n25625), 
         .Z(n41351)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2007[30:82])
    defparam i1_2_lut_rep_264_3_lut.init = 16'h7070;
    FD1P3AX branch_target_m_i2_i25 (.D(branch_target_m_31__N_1157[23]), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(branch_target_m[25])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i25.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_393 (.A(n34433), .B(n39892), .C(n39222), .D(n2_adj_3903), 
         .Z(raw_m_0)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i1_4_lut_adj_393.init = 16'h0002;
    LUT4 operand_w_31__I_0_i5_3_lut (.A(operand_w[4]), .B(multiplier_result_w[4]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i5_3_lut.init = 16'hcaca;
    FD1P3AX branch_target_m_i2_i24 (.D(branch_target_m_31__N_1157[22]), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(branch_target_m[24])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i24.GSR = "ENABLED";
    LUT4 non_debug_exception_w_I_0_2_lut_rep_386 (.A(non_debug_exception_w), 
         .B(valid_w), .Z(n41473)) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2008[34:90])
    defparam non_debug_exception_w_I_0_2_lut_rep_386.init = 16'h8888;
    LUT4 i21141_3_lut_4_lut (.A(non_debug_exception_w), .B(valid_w), .C(ie), 
         .D(operand_1_x[1]), .Z(n23750)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2008[34:90])
    defparam i21141_3_lut_4_lut.init = 16'hf780;
    LUT4 i37811_2_lut (.A(write_idx_m[0]), .B(read_idx_0_d[0]), .Z(n39892)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(470[26:38])
    defparam i37811_2_lut.init = 16'h6666;
    LUT4 m_result_31__I_0_i19_3_lut (.A(m_result[18]), .B(operand_w_31__N_1187[18]), 
         .C(n42746), .Z(operand_w_31__N_840[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i19_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_rep_387 (.A(csr_x[2]), .B(csr_x[4]), .C(csr_x[3]), .Z(n41474)) /* synthesis lut_function=(A+(B+(C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i2_3_lut_rep_387.init = 16'hfefe;
    LUT4 i36671_3_lut (.A(write_idx_m[4]), .B(n39142), .C(read_idx_0_d[4]), 
         .Z(n39222)) /* synthesis lut_function=(A (B+!(C))+!A (B+(C))) */ ;
    defparam i36671_3_lut.init = 16'hdede;
    LUT4 csr_x_0__bdd_2_lut_38190_4_lut (.A(csr_x[2]), .B(csr_x[4]), .C(csr_x[3]), 
         .D(csr_x[1]), .Z(n39068)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam csr_x_0__bdd_2_lut_38190_4_lut.init = 16'hfffe;
    LUT4 mux_19174_i17_3_lut (.A(pc_m[18]), .B(memop_pc_w[18]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i17_3_lut.init = 16'hcaca;
    LUT4 write_idx_m_4__I_0_747_i2_2_lut (.A(write_idx_m[1]), .B(read_idx_0_d[1]), 
         .Z(n2_adj_3903)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1486[18:47])
    defparam write_idx_m_4__I_0_747_i2_2_lut.init = 16'h6666;
    FD1P3AX branch_target_m_i2_i23 (.D(branch_target_m_31__N_1157[21]), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(branch_target_m[23])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i23.GSR = "ENABLED";
    LUT4 operand_w_31__I_0_i10_3_lut (.A(operand_w[9]), .B(multiplier_result_w[9]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i10_3_lut.init = 16'hcaca;
    FD1P3AX branch_target_m_i2_i22 (.D(branch_target_m_31__N_1157[20]), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(branch_target_m[22])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i22.GSR = "ENABLED";
    LUT4 i36595_4_lut (.A(write_idx_m[3]), .B(write_idx_m[2]), .C(read_idx_0_d[3]), 
         .D(read_idx_0_d[2]), .Z(n39142)) /* synthesis lut_function=(!(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D))))) */ ;
    defparam i36595_4_lut.init = 16'h7bde;
    LUT4 mux_20532_i3_3_lut (.A(n23054), .B(n23086), .C(read_idx_0_d[4]), 
         .Z(n23116[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i3_3_lut.init = 16'hcaca;
    LUT4 size_x_1__I_0_153_Mux_30_i3_3_lut_4_lut_4_lut (.A(condition_x[0]), 
         .B(n2_adj_3904), .C(size_x[1]), .D(store_operand_x[6]), .Z(store_data_x[30])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam size_x_1__I_0_153_Mux_30_i3_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 size_x_1__I_0_153_Mux_14_i3_3_lut_4_lut_4_lut (.A(condition_x[0]), 
         .B(store_operand_x[14]), .C(size_x[1]), .D(store_operand_x[6]), 
         .Z(store_data_x[14])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam size_x_1__I_0_153_Mux_14_i3_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 size_x_1__I_0_153_Mux_15_i3_3_lut_4_lut_4_lut (.A(condition_x[0]), 
         .B(store_operand_x[15]), .C(size_x[1]), .D(store_operand_x[7]), 
         .Z(store_data_x[15])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam size_x_1__I_0_153_Mux_15_i3_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 m_result_31__I_0_i32_3_lut (.A(m_result[31]), .B(operand_w_31__N_1187[31]), 
         .C(n42746), .Z(operand_w_31__N_840[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i32_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_394 (.A(n29325), .B(n36706), .C(jrx_csr_read_data[1]), 
         .D(n41432), .Z(csr_read_data_x[1])) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_394.init = 16'hfeee;
    LUT4 mux_19174_i30_3_lut (.A(pc_m[31]), .B(memop_pc_w[31]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i30_3_lut.init = 16'hcaca;
    FD1P3AX branch_target_m_i2_i21 (.D(branch_target_m_31__N_1157[19]), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(branch_target_m[21])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i21.GSR = "ENABLED";
    LUT4 size_x_1__I_0_153_Mux_31_i3_3_lut_4_lut_4_lut (.A(condition_x[0]), 
         .B(n2_adj_3905), .C(size_x[1]), .D(store_operand_x[7]), .Z(store_data_x[31])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam size_x_1__I_0_153_Mux_31_i3_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i1_4_lut_adj_395 (.A(eie), .B(n39068), .C(im[1]), .D(csr_x[0]), 
         .Z(n36706)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_395.init = 16'h3022;
    FD1P3AX condition_met_m_674 (.D(condition_met_x), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(condition_met_m));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam condition_met_m_674.GSR = "ENABLED";
    LUT4 i37221_4_lut_4_lut (.A(condition_x[0]), .B(size_x[1]), .C(n24748), 
         .D(cmp_zero), .Z(n39775)) /* synthesis lut_function=(A (B (C)+!B (D))+!A ((C)+!B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam i37221_4_lut_4_lut.init = 16'hf3d1;
    LUT4 operand_w_31__I_0_i9_3_lut (.A(operand_w[8]), .B(multiplier_result_w[8]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 i37851_2_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), .Z(n39459)) /* synthesis lut_function=(A+(B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1607[18] 1621[32])
    defparam i37851_2_lut.init = 16'heeee;
    FD1P3AX m_result_sel_compare_m_661_rep_449 (.D(m_result_sel_compare_x), 
            .SP(w_clk_cpu_enable_985), .CK(w_clk_cpu), .Q(n42730));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam m_result_sel_compare_m_661_rep_449.GSR = "ENABLED";
    LUT4 m_result_31__I_0_i18_3_lut (.A(m_result[17]), .B(operand_w_31__N_1187[17]), 
         .C(n42746), .Z(operand_w_31__N_840[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i18_3_lut.init = 16'hcaca;
    LUT4 mux_20532_i9_3_lut (.A(n23060), .B(n23092), .C(read_idx_0_d[4]), 
         .Z(n23116[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i9_3_lut.init = 16'hcaca;
    FD1P3AX branch_target_m_i2_i20 (.D(branch_target_m_31__N_1157[18]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(branch_target_m[20])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i20.GSR = "ENABLED";
    LUT4 mux_19174_i16_3_lut (.A(pc_m[17]), .B(memop_pc_w[17]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i16_3_lut.init = 16'hcaca;
    LUT4 mux_20532_i10_3_lut (.A(n23061), .B(n23093), .C(read_idx_0_d[4]), 
         .Z(n23116[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i10_3_lut.init = 16'hcaca;
    LUT4 m_result_31__I_0_i31_3_lut (.A(m_result[30]), .B(operand_w_31__N_1187[30]), 
         .C(n42746), .Z(operand_w_31__N_840[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i31_3_lut.init = 16'hcaca;
    LUT4 mux_19174_i29_3_lut (.A(pc_m[30]), .B(memop_pc_w[30]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i29_3_lut.init = 16'hcaca;
    LUT4 mux_20532_i11_3_lut (.A(n23062), .B(n23094), .C(read_idx_0_d[4]), 
         .Z(n23116[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i11_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_396 (.A(n29325), .B(n36708), .C(jrx_csr_read_data[2]), 
         .D(n41432), .Z(csr_read_data_x[2])) /* synthesis lut_function=(A+(B+(C (D)))) */ ;
    defparam i1_4_lut_adj_396.init = 16'hfeee;
    LUT4 i1_4_lut_adj_397 (.A(bie), .B(n39068), .C(im[2]), .D(csr_x[0]), 
         .Z(n36708)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam i1_4_lut_adj_397.init = 16'h3022;
    LUT4 mux_20532_i12_3_lut (.A(n23063), .B(n23095), .C(read_idx_0_d[4]), 
         .Z(n23116[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i12_3_lut.init = 16'hcaca;
    FD1P3AX branch_target_m_i2_i19 (.D(branch_target_m_31__N_1157[17]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(branch_target_m[19])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i19.GSR = "ENABLED";
    FD1P3AX m_result_sel_compare_m_661 (.D(m_result_sel_compare_x), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(m_result_sel_compare_m));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam m_result_sel_compare_m_661.GSR = "ENABLED";
    LUT4 mux_20532_i13_3_lut (.A(n23064), .B(n23096), .C(read_idx_0_d[4]), 
         .Z(n23116[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i13_3_lut.init = 16'hcaca;
    LUT4 m_result_31__I_0_i30_3_lut (.A(m_result[29]), .B(operand_w_31__N_1187[29]), 
         .C(n42746), .Z(operand_w_31__N_840[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i30_3_lut.init = 16'hcaca;
    LUT4 mux_19174_i28_3_lut (.A(pc_m[29]), .B(memop_pc_w[29]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i28_3_lut.init = 16'hcaca;
    LUT4 mux_20532_i14_3_lut (.A(n23065), .B(n23097), .C(read_idx_0_d[4]), 
         .Z(n23116[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i14_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i8_3_lut (.A(operand_w[7]), .B(multiplier_result_w[7]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i4_3_lut (.A(operand_w[3]), .B(multiplier_result_w[3]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 m_result_31__I_0_i29_3_lut (.A(m_result[28]), .B(operand_w_31__N_1187[28]), 
         .C(n42746), .Z(operand_w_31__N_840[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i29_3_lut.init = 16'hcaca;
    LUT4 mux_19174_i27_3_lut (.A(pc_m[28]), .B(memop_pc_w[28]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i27_3_lut.init = 16'hcaca;
    FD1P3AX branch_target_m_i2_i18 (.D(branch_target_m_31__N_1157[16]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(branch_target_m[18])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i18.GSR = "ENABLED";
    FD1P3AX branch_target_m_i2_i17 (.D(branch_target_m_31__N_1157[15]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(branch_target_m[17])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i17.GSR = "ENABLED";
    LUT4 mux_20532_i15_3_lut (.A(n23066), .B(n23098), .C(read_idx_0_d[4]), 
         .Z(n23116[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i15_3_lut.init = 16'hcaca;
    LUT4 mux_20532_i1_3_lut (.A(n23052), .B(n23084), .C(read_idx_0_d[4]), 
         .Z(n23116[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i1_3_lut.init = 16'hcaca;
    LUT4 mux_75_i26_3_lut (.A(logic_result_x[25]), .B(mc_result_x[25]), 
         .C(x_result_sel_mc_arith_x), .Z(n1253[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1619[18] 1621[32])
    defparam mux_75_i26_3_lut.init = 16'hcaca;
    FD1P3AX branch_target_m_i2_i16 (.D(branch_target_m_31__N_1157[14]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(branch_target_m[16])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i16.GSR = "ENABLED";
    LUT4 m_result_31__I_0_i28_3_lut (.A(m_result[27]), .B(operand_w_31__N_1187[27]), 
         .C(n42746), .Z(operand_w_31__N_840[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i28_3_lut.init = 16'hcaca;
    LUT4 mux_19174_i26_3_lut (.A(pc_m[27]), .B(memop_pc_w[27]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i26_3_lut.init = 16'hcaca;
    LUT4 mux_20532_i4_3_lut (.A(n23055), .B(n23087), .C(read_idx_0_d[4]), 
         .Z(n23116[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i4_3_lut.init = 16'hcaca;
    LUT4 i22_4_lut_3_lut (.A(csr_x[0]), .B(jrx_csr_read_data[0]), .C(csr_x[3]), 
         .Z(n9)) /* synthesis lut_function=(A (B (C))+!A !(C)) */ ;
    defparam i22_4_lut_3_lut.init = 16'h8585;
    LUT4 i2_3_lut_4_lut_4_lut (.A(csr_x[0]), .B(n31712), .C(n41391), .D(csr_write_enable_x), 
         .Z(dc_re_N_2934)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2_3_lut_4_lut_4_lut.init = 16'h1000;
    LUT4 i1_2_lut_3_lut_3_lut (.A(csr_x[0]), .B(n41503), .C(csr_x[3]), 
         .Z(n29325)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i1_2_lut_3_lut_3_lut.init = 16'h0404;
    LUT4 i1_3_lut_4_lut_4_lut (.A(csr_x[0]), .B(eba[11]), .C(csr_x[1]), 
         .D(csr_x[3]), .Z(n30)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((D)+!C))) */ ;
    defparam i1_3_lut_4_lut_4_lut.init = 16'h00d0;
    LUT4 i1_2_lut_4_lut_adj_398 (.A(csr_x[1]), .B(csr_x[3]), .C(csr_x[0]), 
         .D(deba[11]), .Z(n29)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_2_lut_4_lut_adj_398.init = 16'h4000;
    FD1P3AX branch_target_m_i2_i15 (.D(branch_target_m_31__N_1157[13]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(branch_target_m[15])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i15.GSR = "ENABLED";
    FD1P3AX branch_target_m_i2_i14 (.D(branch_target_m_31__N_1157[12]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(branch_target_m[14])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i14.GSR = "ENABLED";
    LUT4 m_result_31__I_0_i27_3_lut (.A(m_result[26]), .B(operand_w_31__N_1187[26]), 
         .C(n42746), .Z(operand_w_31__N_840[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i27_3_lut.init = 16'hcaca;
    LUT4 mux_19174_i25_3_lut (.A(pc_m[26]), .B(memop_pc_w[26]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i25_3_lut.init = 16'hcaca;
    LUT4 operand_w_31__I_0_i7_3_lut (.A(operand_w[6]), .B(multiplier_result_w[6]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i7_3_lut.init = 16'hcaca;
    LUT4 mux_20532_i26_3_lut (.A(n23077), .B(n23109), .C(read_idx_0_d[4]), 
         .Z(n23116[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i26_3_lut.init = 16'hcaca;
    LUT4 m_result_31__I_0_i26_3_lut (.A(m_result[25]), .B(operand_w_31__N_1187[25]), 
         .C(n42746), .Z(operand_w_31__N_840[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i26_3_lut.init = 16'hcaca;
    LUT4 mux_19174_i24_3_lut (.A(pc_m[25]), .B(memop_pc_w[25]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i24_3_lut.init = 16'hcaca;
    FD1P3AX branch_target_m_i2_i13 (.D(branch_target_m_31__N_1157[11]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(branch_target_m[13])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i13.GSR = "ENABLED";
    FD1P3AX break_x_652 (.D(break_d), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(break_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam break_x_652.GSR = "ENABLED";
    LUT4 mux_20532_i27_3_lut (.A(n23078), .B(n23110), .C(read_idx_0_d[4]), 
         .Z(n23116[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i27_3_lut.init = 16'hcaca;
    LUT4 mux_20532_i28_3_lut (.A(n23079), .B(n23111), .C(read_idx_0_d[4]), 
         .Z(n23116[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i28_3_lut.init = 16'hcaca;
    LUT4 mux_20532_i29_3_lut (.A(n23080), .B(n23112), .C(read_idx_0_d[4]), 
         .Z(n23116[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i29_3_lut.init = 16'hcaca;
    LUT4 m_result_31__I_0_i25_3_lut (.A(m_result[24]), .B(operand_w_31__N_1187[24]), 
         .C(n42746), .Z(operand_w_31__N_840[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i25_3_lut.init = 16'hcaca;
    LUT4 mux_19174_i23_3_lut (.A(pc_m[24]), .B(memop_pc_w[24]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i23_3_lut.init = 16'hcaca;
    FD1P3AX branch_target_m_i2_i12 (.D(branch_target_m_31__N_1157[10]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(branch_target_m[12])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i12.GSR = "ENABLED";
    FD1P3AX branch_target_m_i2_i11 (.D(branch_target_m_31__N_1157[9]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(branch_target_m[11])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i11.GSR = "ENABLED";
    LUT4 mux_20532_i30_3_lut (.A(n23081), .B(n23113), .C(read_idx_0_d[4]), 
         .Z(n23116[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i30_3_lut.init = 16'hcaca;
    FD1P3AX direction_x_647 (.D(logic_op_d[3]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(direction_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam direction_x_647.GSR = "ENABLED";
    LUT4 mux_20532_i31_3_lut (.A(n23082), .B(n23114), .C(read_idx_0_d[4]), 
         .Z(n23116[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i31_3_lut.init = 16'hcaca;
    LUT4 mux_20532_i32_3_lut (.A(n23083), .B(n23115), .C(read_idx_0_d[4]), 
         .Z(n23116[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_20532_i32_3_lut.init = 16'hcaca;
    LUT4 m_result_31__I_0_i24_3_lut (.A(m_result[23]), .B(operand_w_31__N_1187[23]), 
         .C(n42746), .Z(operand_w_31__N_840[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i24_3_lut.init = 16'hcaca;
    FD1P3AX branch_target_m_i2_i10 (.D(branch_target_m_31__N_1157[8]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(branch_target_m[10])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i10.GSR = "ENABLED";
    FD1P3AX branch_target_m_i2_i9 (.D(branch_target_m_31__N_1157[7]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(branch_target_m[9])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i9.GSR = "ENABLED";
    FD1P3AX branch_target_m_i2_i8 (.D(branch_target_m_31__N_1157[6]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(branch_target_m[8])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i8.GSR = "ENABLED";
    LUT4 mux_19174_i22_3_lut (.A(pc_m[23]), .B(memop_pc_w[23]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i22_3_lut.init = 16'hcaca;
    LUT4 m_result_31__I_0_i23_3_lut (.A(m_result[22]), .B(operand_w_31__N_1187[22]), 
         .C(n42746), .Z(operand_w_31__N_840[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i23_3_lut.init = 16'hcaca;
    LUT4 mux_19174_i21_3_lut (.A(pc_m[22]), .B(memop_pc_w[22]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i21_3_lut.init = 16'hcaca;
    PFUMX i38 (.BLUT(n29), .ALUT(n30), .C0(csr_x[2]), .Z(n31));
    LUT4 m_result_31__I_0_i22_3_lut (.A(m_result[21]), .B(operand_w_31__N_1187[21]), 
         .C(n42746), .Z(operand_w_31__N_840[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i22_3_lut.init = 16'hcaca;
    PFUMX i38619 (.BLUT(n41612), .ALUT(n41613), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[21]));
    LUT4 mux_19174_i20_3_lut (.A(pc_m[21]), .B(memop_pc_w[21]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i20_3_lut.init = 16'hcaca;
    PFUMX i38617 (.BLUT(n41609), .ALUT(n41610), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[28]));
    FD1P3AX branch_target_m_i2_i7 (.D(branch_target_m_31__N_1157[5]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(branch_target_m[7])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i7.GSR = "ENABLED";
    FD1P3AX sign_extend_x_643 (.D(instruction[28]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(sign_extend_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam sign_extend_x_643.GSR = "ENABLED";
    PFUMX i38615 (.BLUT(n41606), .ALUT(n41607), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[16]));
    LUT4 m_result_31__I_0_i21_3_lut (.A(m_result[20]), .B(operand_w_31__N_1187[20]), 
         .C(n42746), .Z(operand_w_31__N_840[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[25:125])
    defparam m_result_31__I_0_i21_3_lut.init = 16'hcaca;
    PFUMX i38613 (.BLUT(n41603), .ALUT(n41604), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[17]));
    LUT4 mux_19174_i19_3_lut (.A(pc_m[20]), .B(memop_pc_w[20]), .C(data_bus_error_exception_m), 
         .Z(operand_w_31__N_1187[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2594[48:114])
    defparam mux_19174_i19_3_lut.init = 16'hcaca;
    PFUMX i38611 (.BLUT(n41600), .ALUT(n41601), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[27]));
    PFUMX i38609 (.BLUT(n41597), .ALUT(n41598), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[26]));
    LUT4 i29225_3_lut_4_lut (.A(bus_error_x), .B(valid_x), .C(n41526), 
         .D(data_bus_error_exception), .Z(eid_x_2__N_999[2])) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A ((D)+!C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1750[42] 1752[43])
    defparam i29225_3_lut_4_lut.init = 16'hff07;
    PFUMX i38607 (.BLUT(n41594), .ALUT(n41595), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[25]));
    PFUMX i38605 (.BLUT(n41591), .ALUT(n41592), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[24]));
    FD1P3AX branch_target_m_i2_i6 (.D(branch_target_m_31__N_1157[4]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(branch_target_m[6])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i6.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut_adj_399 (.A(bus_error_x), .B(valid_x), .C(n41526), 
         .D(divide_by_zero_x), .Z(n38801)) /* synthesis lut_function=(!(A (B (C)+!B (C+(D)))+!A (C+(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1750[42] 1752[43])
    defparam i1_3_lut_4_lut_adj_399.init = 16'h080f;
    FD1P3AX branch_target_m_i2_i5 (.D(branch_target_m_31__N_1157[3]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(branch_target_m[5])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam branch_target_m_i2_i5.GSR = "ENABLED";
    PFUMX i38603 (.BLUT(n41588), .ALUT(n41589), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[23]));
    FD1P3AX load_x_640 (.D(n41384), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(load_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam load_x_640.GSR = "ENABLED";
    PFUMX i38601 (.BLUT(n41585), .ALUT(n41586), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[22]));
    PFUMX i38599 (.BLUT(n41582), .ALUT(n41583), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[20]));
    LUT4 operand_w_31__I_0_i6_3_lut (.A(operand_w[5]), .B(multiplier_result_w[5]), 
         .C(w_result_sel_mul_w), .Z(w_result_31__N_680[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1639[19] 1641[28])
    defparam operand_w_31__I_0_i6_3_lut.init = 16'hcaca;
    PFUMX i38597 (.BLUT(n41579), .ALUT(n41580), .C0(non_debug_exception_x_N_1357), 
          .Z(branch_target_m_31__N_1157[19]));
    FD1P3AX x_result_sel_csr_x_626 (.D(x_result_sel_csr_d), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(x_result_sel_csr_x));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam x_result_sel_csr_x_626.GSR = "ENABLED";
    FD1P3AX csr_x_i0_i4 (.D(read_idx_0_d[4]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(csr_x[4])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam csr_x_i0_i4.GSR = "ENABLED";
    FD1P3AX csr_x_i0_i3 (.D(read_idx_0_d[3]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(csr_x[3])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam csr_x_i0_i3.GSR = "ENABLED";
    FD1P3AX csr_x_i0_i2 (.D(read_idx_0_d[2]), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(csr_x[2])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2418[5] 2626[8])
    defparam csr_x_i0_i2.GSR = "ENABLED";
    PFUMX i23_adj_400 (.BLUT(n3_adj_3816), .ALUT(n7_adj_3796), .C0(csr_x[3]), 
          .Z(n10_adj_3897));
    PFUMX m_result_31__I_0_705_i1 (.BLUT(shifter_result_m[0]), .ALUT(m_result_31__N_648[0]), 
          .C0(n39334), .Z(m_result[0])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    CCU2D operand_0_x_31__I_0_0 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(operand_1_x[31]), .B1(muliplicand[31]), .C1(operand_1_x[30]), 
          .D1(muliplicand[30]), .COUT(n36486));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1585[19:45])
    defparam operand_0_x_31__I_0_0.INIT0 = 16'hF000;
    defparam operand_0_x_31__I_0_0.INIT1 = 16'h9009;
    defparam operand_0_x_31__I_0_0.INJECT1_0 = "NO";
    defparam operand_0_x_31__I_0_0.INJECT1_1 = "YES";
    PFUMX w_result_31__I_0_i2 (.BLUT(w_result_31__N_680[1]), .ALUT(load_data_w[1]), 
          .C0(w_result_sel_load_w), .Z(w_result[1])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=10, LSE_RCOL=6, LSE_LLINE=283, LSE_RLINE=366 */ ;
    lm32_shifter shifter (.left_shift_result({left_shift_result}), .w_clk_cpu(w_clk_cpu), 
            .w_clk_cpu_enable_984(w_clk_cpu_enable_984), .\operand_1_x[4] (operand_1_x[4]), 
            .\operand_1_x[2] (operand_1_x[2]), .\operand_1_x[3] (operand_1_x[3]), 
            .direction_m(direction_m), .shifter_result_m({shifter_result_m}), 
            .\operand_1_x[1] (operand_1_x[1]), .\operand_1_x[0] (operand_1_x[0]), 
            .muliplicand({muliplicand}), .direction_x(direction_x), .sign_extend_x(sign_extend_x)) /* synthesis syn_module_defined=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1071[14] 1082[6])
    lm32_multiplier multiplier (.GND_net(GND_net), .muliplicand({muliplicand}), 
            .operand_1_x({operand_1_x}), .multiplier_result_w({multiplier_result_w}), 
            .w_clk_cpu(w_clk_cpu), .n41428(n41428), .store_m(store_m), 
            .LM32D_CYC_O(LM32D_CYC_O), .n41512(n41512), .w_clk_cpu_enable_623(w_clk_cpu_enable_623), 
            .n46(n46), .reset_exception(reset_exception), .n22524(n22524), 
            .\size_x[1] (size_x[1]), .\condition_x[0] (condition_x[0]), 
            .n26122(n26122), .n41513(n41513), .data_bus_error_exception(data_bus_error_exception), 
            .memop_pc_w_31__N_1219(memop_pc_w_31__N_1219), .w_clk_cpu_enable_972(w_clk_cpu_enable_972), 
            .w_clk_cpu_enable_984(w_clk_cpu_enable_984), .n26142(n26142), 
            .\bypass_data_0[1] (bypass_data_0[1]), .w_clk_cpu_enable_711(w_clk_cpu_enable_711), 
            .\bypass_data_0[0] (bypass_data_0[0]), .\d_result_0[31] (d_result_0[31]), 
            .\d_result_0[30] (d_result_0[30]), .\d_result_0[29] (d_result_0[29]), 
            .\d_result_0[28] (d_result_0[28]), .\d_result_0[27] (d_result_0[27]), 
            .\d_result_0[26] (d_result_0[26]), .\d_result_0[25] (d_result_0[25]), 
            .\d_result_0[24] (d_result_0[24]), .\d_result_0[23] (d_result_0[23]), 
            .\d_result_0[22] (d_result_0[22]), .\d_result_0[21] (d_result_0[21]), 
            .\d_result_0[20] (d_result_0[20]), .\d_result_0[19] (d_result_0[19]), 
            .\d_result_0[18] (d_result_0[18]), .\d_result_0[17] (d_result_0[17]), 
            .\d_result_0[16] (d_result_0[16]), .\d_result_0[15] (d_result_0[15]), 
            .\d_result_0[14] (d_result_0[14]), .\d_result_0[13] (d_result_0[13]), 
            .\d_result_0[12] (d_result_0[12]), .\d_result_0[11] (d_result_0[11]), 
            .\d_result_0[10] (d_result_0[10]), .\d_result_0[9] (d_result_0[9]), 
            .\d_result_0[8] (d_result_0[8]), .\d_result_0[7] (d_result_0[7]), 
            .\d_result_0[6] (d_result_0[6]), .\d_result_0[5] (d_result_0[5]), 
            .\d_result_0[4] (d_result_0[4]), .\d_result_0[3] (d_result_0[3]), 
            .\d_result_0[2] (d_result_0[2])) /* synthesis syn_module_defined=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1087[17] 1097[6])
    lm32_mc_arithmetic mc_arithmetic (.reg_data_1({reg_data_1}), .w_result({w_result}), 
            .n18863(n18863), .operand_m({operand_m}), .left_shift_result({left_shift_result}), 
            .m_result_sel_shift_m(m_result_sel_shift_m), .n1826({n1826[31:24], 
            Open_38, Open_39, Open_40, Open_41, Open_42, Open_43, 
            Open_44, Open_45, Open_46, Open_47, Open_48, Open_49, 
            Open_50, n1826[10:8], Open_51, Open_52, Open_53, Open_54, 
            Open_55, Open_56, Open_57, Open_58}), .n18875(n18875), 
            .w_clk_cpu(w_clk_cpu), .w_clk_cpu_enable_958(w_clk_cpu_enable_958), 
            .n41406(n41406), .n37259(n37259), .n41391(n41391), .load_x(load_x), 
            .n39970(n39970), .bypass_data_0({bypass_data_0}), .n41417(n41417), 
            .w_clk_cpu_enable_865(w_clk_cpu_enable_865), .mc_result_x({mc_result_x}), 
            .mc_stall_request_x(mc_stall_request_x), .GND_net(GND_net), 
            .n21435(n21411[0]), .n21434(n21411[1]), .n21433(n21411[2]), 
            .n21432(n21411[3]), .n21431(n21411[4]), .n21430(n21411[5]), 
            .n21429(n21411[6]), .n1857(n1826[1]), .n1856(n1826[2]), .n1855(n1826[3]), 
            .n1854(n1826[4]), .n1853(n1826[5]), .n41364(n41364), .n22236(n22236), 
            .\instruction_d[11] (instruction_d[11]), .n41380(n41380), .n2(n2_adj_3889), 
            .n1852(n1826[6]), .n18869(n18869), .\instruction_d[12] (instruction_d[12]), 
            .n2_adj_50(n2_adj_3887), .n1851(n1826[7]), .\instruction_d[13] (instruction_d[13]), 
            .n2_adj_51(n2_adj_3885), .\instruction_d[14] (instruction_d[14]), 
            .n2_adj_52(n2_adj_3883), .sign_extend_immediate(sign_extend_immediate), 
            .\instruction_d[15] (instruction_d[15]), .n36772(n36772), .\instruction_d[0] (instruction_d[0]), 
            .n2_adj_53(n2_adj_3840), .\instruction_d[1] (instruction_d[1]), 
            .n2_adj_54(n2_adj_3838), .\instruction_d[2] (instruction_d[2]), 
            .n2_adj_55(n2_adj_3836), .\instruction_d[3] (instruction_d[3]), 
            .n2_adj_56(n2_adj_3833), .\instruction_d[4] (instruction_d[4]), 
            .n2_adj_57(n2_adj_3831), .\instruction_d[5] (instruction_d[5]), 
            .n2_adj_58(n2_adj_3829), .\instruction_d[6] (instruction_d[6]), 
            .n2_adj_59(n2_adj_3827), .\instruction_d[7] (instruction_d[7]), 
            .n2_adj_60(n2_adj_3825), .\instruction_d[8] (instruction_d[8]), 
            .n2_adj_61(n2_adj_3823), .\instruction_d[9] (instruction_d[9]), 
            .n2_adj_62(n2_adj_3821), .\instruction_d[10] (instruction_d[10]), 
            .n2_adj_63(n2), .divide_by_zero_x(divide_by_zero_x), .condition_met_m(condition_met_m), 
            .m_result_sel_compare_m(m_result_sel_compare_m), .n41367(n41367), 
            .raw_x_1(raw_x_1), .cycles_5__N_2495(cycles_5__N_2495), .csr_read_data_x({csr_read_data_x}), 
            .adder_result_x({adder_result_x}), .x_result_sel_add_x(x_result_sel_add_x), 
            .\x_result_31__N_616[1] (x_result_31__N_616[1]), .\x_result_31__N_616[2] (x_result_31__N_616[2]), 
            .\x_result_31__N_616[3] (x_result_31__N_616[3]), .\x_result_31__N_616[4] (x_result_31__N_616[4]), 
            .\x_result_31__N_616[5] (x_result_31__N_616[5]), .\x_result_31__N_616[6] (x_result_31__N_616[6]), 
            .\x_result_31__N_616[7] (x_result_31__N_616[7]), .\x_result_31__N_616[15] (x_result_31__N_616[15]), 
            .n13(n13), .\x_result_31__N_616[16] (x_result_31__N_616[16]), 
            .\x_result_31__N_616[17] (x_result_31__N_616[17]), .n41373(n41373), 
            .n41408(n41408), .\x_result_31__N_616[18] (x_result_31__N_616[18]), 
            .\x_result_31__N_616[19] (x_result_31__N_616[19]), .\x_result_31__N_616[20] (x_result_31__N_616[20]), 
            .\x_result_31__N_616[21] (x_result_31__N_616[21]), .\x_result_31__N_616[22] (x_result_31__N_616[22]), 
            .x_result_sel_csr_x(x_result_sel_csr_x), .x_result_sel_sext_x(x_result_sel_sext_x), 
            .n41411(n41411), .direction_m(direction_m), .n41407(n41407), 
            .pc_f({pc_f}), .\x_result_31__N_616[23] (x_result_31__N_616[23]), 
            .\x_result_31__N_616[24] (x_result_31__N_616[24]), .\x_result_31__N_616[25] (x_result_31__N_616[25]), 
            .n42740(n42740), .n41361(n41361), .\x_result_31__N_616[26] (x_result_31__N_616[26]), 
            .\x_result_31__N_616[27] (x_result_31__N_616[27]), .\x_result_31__N_616[28] (x_result_31__N_616[28]), 
            .\x_result_31__N_616[0] (x_result_31__N_616[0]), .\x_result_31__N_616[29] (x_result_31__N_616[29]), 
            .\x_result_31__N_616[30] (x_result_31__N_616[30]), .\x_result_31__N_616[31] (x_result_31__N_616[31]), 
            .w_clk_cpu_enable_984(w_clk_cpu_enable_984), .LM32I_CYC_O(LM32I_CYC_O), 
            .i_cyc_o_N_1759(i_cyc_o_N_1759), .w_clk_cpu_enable_216(w_clk_cpu_enable_216), 
            .n21414(n21411[21]), .n37179(n37179), .\muliplicand[0] (muliplicand[0]), 
            .n1285(n1253[0]), .\muliplicand[7] (muliplicand[7]), .\muliplicand[6] (muliplicand[6]), 
            .\muliplicand[5] (muliplicand[5]), .\muliplicand[4] (muliplicand[4]), 
            .\muliplicand[3] (muliplicand[3]), .n41345(n41345), .\muliplicand[2] (muliplicand[2]), 
            .\muliplicand[1] (muliplicand[1]), .n1844(n1826[14]), .n1845(n1826[13]), 
            .n1846(n1826[12]), .n1847(n1826[11]), .n38799(n38799), .n38840(n38840), 
            .n1791(n1760[1]), .n1790(n1760[2]), .n1789(n1760[3]), .n1788(n1760[4]), 
            .n1787(n1760[5]), .n1786(n1760[6]), .n1785(n1760[7]), .n1777(n1760[15]), 
            .n1776(n1760[16]), .n1775(n1760[17]), .n1774(n1760[18]), .n1773(n1760[19]), 
            .n1772(n1760[20]), .n1771(n1760[21]), .n1770(n1760[22]), .n1769(n1760[23]), 
            .n1768(n1760[24]), .n1767(n1760[25]), .n1766(n1760[26]), .n1765(n1760[27]), 
            .n1764(n1760[28]), .n1792(n1760[0]), .n1763(n1760[29]), .n1762(n1760[30]), 
            .n1843(n1826[15]), .n1842(n1826[16]), .n1841(n1826[17]), .n1840(n1826[18]), 
            .n1839(n1826[19]), .n1838(n1826[20]), .n1837(n1826[21]), .n1836(n1826[22]), 
            .n1835(n1826[23])) /* synthesis syn_module_defined=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1102[20] 1128[6])
    lm32_logic_op logic_op (.\logic_op_x[2] (logic_op_x[2]), .\logic_op_x[3] (logic_op_x[3]), 
            .muliplicand({muliplicand}), .\condition_x[0] (condition_x[0]), 
            .\size_x[1] (size_x[1]), .operand_1_x({operand_1_x}), .logic_result_x({logic_result_x})) /* synthesis syn_module_defined=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1059[15] 1067[6])
    lm32_load_store_unit load_store_unit (.store_operand_x({store_operand_x}), 
            .\condition_x[0] (condition_x[0]), .\size_x[1] (size_x[1]), 
            .wb_load_complete(wb_load_complete), .w_clk_cpu(w_clk_cpu), 
            .w_clk_cpu_enable_972(w_clk_cpu_enable_972), .LM32D_WE_O(LM32D_WE_O), 
            .w_clk_cpu_enable_886(w_clk_cpu_enable_886), .n41372(n41372), 
            .LM32D_DAT_O({LM32D_DAT_O}), .w_clk_cpu_enable_623(w_clk_cpu_enable_623), 
            .SHAREDBUS_DAT_O({SHAREDBUS_DAT_O}), .LM32D_ADR_O({LM32D_ADR_O}), 
            .operand_m({operand_m}), .LM32D_SEL_O({LM32D_SEL_O}), .LM32D_STB_O(LM32D_STB_O), 
            .w_clk_cpu_enable_245(w_clk_cpu_enable_245), .n41492(n41492), 
            .byte_enable_x({Open_59, Open_60, Open_61, byte_enable_x[0]}), 
            .LM32D_CYC_O(LM32D_CYC_O), .n26096(n26096), .n26122(n26122), 
            .\operand_w[0] (operand_w[0]), .load_data_w({load_data_w}), 
            .\operand_w[1] (operand_w[1]), .n2(n2_adj_3905), .n2_adj_49(n2_adj_3904), 
            .\byte_enable_x[1] (byte_enable_x[1]), .wb_load_complete_N_2129(wb_load_complete_N_2129), 
            .w_clk_cpu_enable_711(w_clk_cpu_enable_711), .stall_wb_load_N_2112(stall_wb_load_N_2112), 
            .n42746(n42746), .n46(n46), .n4(n4_adj_3899), .n41428(n41428), 
            .n41491(n41491), .\adder_result_x[1] (adder_result_x[1]), .\adder_result_x[0] (adder_result_x[0]), 
            .wb_select_m(wb_select_m), .w_clk_cpu_enable_878(w_clk_cpu_enable_878), 
            .n42726(n42726), .\store_data_x[31] (store_data_x[31]), .\store_data_x[30] (store_data_x[30]), 
            .sign_extend_x(sign_extend_x), .w_clk_cpu_enable_985(w_clk_cpu_enable_985), 
            .\store_data_x[15] (store_data_x[15]), .stall_wb_load(stall_wb_load), 
            .exception_m(exception_m), .\store_data_x[14] (store_data_x[14])) /* synthesis syn_module_defined=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(984[5] 1043[6])
    lm32_jtag jtag_reg_d_7__I_0 (.jtag_reg_d({jtag_reg_d}), .w_clk_cpu(w_clk_cpu), 
            .GND_net(GND_net), .n41428(n41428), .n39970(n39970), .branch_flushX_m_N_1116(branch_flushX_m_N_1116), 
            .cycles_5__N_2495(cycles_5__N_2495), .n42740(n42740), .w_clk_cpu_enable_914(w_clk_cpu_enable_914), 
            .n41391(n41391), .load_x(load_x), .n41395(n41395), .stall_wb_load_N_2112(stall_wb_load_N_2112), 
            .w_clk_cpu_enable_697(w_clk_cpu_enable_697), .n26126(n26126), 
            .csr_write_enable_x(csr_write_enable_x), .n41357(n41357), .LM32I_CYC_O(LM32I_CYC_O), 
            .w_clk_cpu_enable_763(w_clk_cpu_enable_763), .branch_taken_m(branch_taken_m), 
            .w_clk_cpu_enable_638(w_clk_cpu_enable_638), .w_clk_cpu_enable_984(w_clk_cpu_enable_984), 
            .n41365(n41365), .\csr_x[0] (csr_x[0]), .n41444(n41444), .n41457(n41457), 
            .eba_31__N_1101(eba_31__N_1101), .\operand_1_x[0] (operand_1_x[0]), 
            .n31712(n31712), .deba_31__N_1120(deba_31__N_1120), .jtag_break(jtag_break), 
            .reset_exception(reset_exception), .\jrx_csr_read_data[0] (jrx_csr_read_data[0]), 
            .jtag_reg_q({jtag_reg_q}), .jtag_update_N_2932(jtag_update_N_2932), 
            .\jtag_reg_addr_d[1] (\jtag_reg_addr_d[1] ), .\jtag_reg_addr_d[0] (\jtag_reg_addr_d[0] ), 
            .w_clk_cpu_enable_330(w_clk_cpu_enable_330), .n42726(n42726), 
            .\jrx_csr_read_data[7] (jrx_csr_read_data[7]), .\jrx_csr_read_data[6] (jrx_csr_read_data[6]), 
            .\jrx_csr_read_data[5] (jrx_csr_read_data[5]), .\jrx_csr_read_data[4] (jrx_csr_read_data[4]), 
            .\jrx_csr_read_data[3] (jrx_csr_read_data[3]), .\jrx_csr_read_data[2] (jrx_csr_read_data[2]), 
            .\jrx_csr_read_data[1] (jrx_csr_read_data[1]), .w_clk_cpu_enable_865(w_clk_cpu_enable_865), 
            .w_clk_cpu_enable_958(w_clk_cpu_enable_958), .x_result_sel_csr_d(x_result_sel_csr_d), 
            .n22501(n22501), .n41417(n41417), .n26142(n26142), .w_clk_cpu_enable_983(w_clk_cpu_enable_983), 
            .jtag_reg_addr_q({jtag_reg_addr_q}), .n38725(n38725), .jtag_reg_d_7__N_505(jtag_reg_d_7__N_505), 
            .\operand_1_x[7] (operand_1_x[7]), .\operand_1_x[6] (operand_1_x[6]), 
            .\operand_1_x[5] (operand_1_x[5]), .\operand_1_x[4] (operand_1_x[4]), 
            .\operand_1_x[3] (operand_1_x[3]), .\operand_1_x[2] (operand_1_x[2]), 
            .\operand_1_x[1] (operand_1_x[1])) /* synthesis syn_module_defined=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1163[11] 1208[6])
    lm32_interrupt interrupt (.im({Open_62, Open_63, Open_64, Open_65, 
            Open_66, Open_67, Open_68, Open_69, Open_70, Open_71, 
            im[21:19], Open_72, Open_73, Open_74, Open_75, Open_76, 
            Open_77, Open_78, Open_79, Open_80, Open_81, Open_82, 
            Open_83, Open_84, Open_85, Open_86, Open_87, Open_88, 
            Open_89, Open_90}), .w_clk_cpu(w_clk_cpu), .operand_1_x({operand_1_x}), 
            .\im[18] (im[18]), .\im[17] (im[17]), .\im[16] (im[16]), .\im[15] (im[15]), 
            .\im[14] (im[14]), .\im[13] (im[13]), .\im[12] (im[12]), .\im[11] (im[11]), 
            .\im[10] (im[10]), .\im[9] (im[9]), .\im[31] (im[31]), .\im[8] (im[8]), 
            .\im[30] (im[30]), .\im[7] (im[7]), .\im[29] (im[29]), .\im[6] (im[6]), 
            .\im[28] (im[28]), .\im[5] (im[5]), .bie(bie), .bie_N_2835(bie_N_2835), 
            .\im[27] (im[27]), .\im[4] (im[4]), .eie(eie), .n23750(n23750), 
            .ie(ie), .\csr_x[0] (csr_x[0]), .n21263(n21231[0]), .\im[26] (im[26]), 
            .\im[3] (im[3]), .n41474(n41474), .\csr_x[1] (csr_x[1]), .n25705(n25705), 
            .\im[25] (im[25]), .\im[2] (im[2]), .\im[24] (im[24]), .\im[1] (im[1]), 
            .\im[23] (im[23]), .n41473(n41473), .n41472(n41472), .n25625(n25625), 
            .bret_q_x(bret_q_x), .w_clk_cpu_enable_984(w_clk_cpu_enable_984), 
            .n4(n4_adj_3898), .jtag_reg_d_7__N_505(jtag_reg_d_7__N_505), 
            .n41359(n41359), .ie_N_2822(ie_N_2822), .n41357(n41357), .n41502(n41502), 
            .\csr_x[2] (csr_x[2]), .n38725(n38725), .\im[22] (im[22]), 
            .w_clk_cpu_enable_330(w_clk_cpu_enable_330), .n41391(n41391), 
            .eret_x(eret_x), .bret_x(bret_x), .n41351(n41351), .ie_N_2821(ie_N_2821)) /* synthesis syn_module_defined=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1133[16] 1158[6])
    lm32_instruction_unit instruction_unit (.pc_d({pc_d}), .w_clk_cpu(w_clk_cpu), 
            .w_clk_cpu_enable_983(w_clk_cpu_enable_983), .pc_f({pc_f}), 
            .\instruction_d[13] (instruction_d[13]), .w_clk_cpu_enable_984(w_clk_cpu_enable_984), 
            .branch_taken_m(branch_taken_m), .w_clk_cpu_enable_914(w_clk_cpu_enable_914), 
            .\instruction_d[12] (instruction_d[12]), .\instruction_d[11] (instruction_d[11]), 
            .\instruction_d[10] (instruction_d[10]), .\instruction_d[9] (instruction_d[9]), 
            .\instruction_d[8] (instruction_d[8]), .\instruction_d[7] (instruction_d[7]), 
            .\instruction_d[6] (instruction_d[6]), .\instruction_d[5] (instruction_d[5]), 
            .\instruction_d[4] (instruction_d[4]), .\instruction_d[3] (instruction_d[3]), 
            .\instruction_d[2] (instruction_d[2]), .GND_net(GND_net), .pc_m({pc_m}), 
            .w_clk_cpu_enable_972(w_clk_cpu_enable_972), .\LM32I_ADR_O[2] (\LM32I_ADR_O[2] ), 
            .w_clk_cpu_enable_763(w_clk_cpu_enable_763), .SHAREDBUS_DAT_O({SHAREDBUS_DAT_O}), 
            .LM32I_CYC_O(LM32I_CYC_O), .n37179(n37179), .\instruction_d[0] (instruction_d[0]), 
            .\selected_1__N_344[0] (\selected_1__N_344[0] ), .w_clk_cpu_enable_216(w_clk_cpu_enable_216), 
            .\instruction_d[1] (instruction_d[1]), .n41375(n41375), .n41504(n41504), 
            .\branch_target_d[3] (branch_target_d[3]), .n42746(n42746), 
            .n41459(n41459), .branch_target_m({branch_target_m}), .i_cyc_o_N_1759(i_cyc_o_N_1759), 
            .valid_d(valid_d), .n41394(n41394), .\LM32I_ADR_O[31] (\LM32I_ADR_O[31] ), 
            .bus_error_f_N_1764(bus_error_f_N_1764), .\LM32I_ADR_O[30] (\LM32I_ADR_O[30] ), 
            .\branch_target_d[30] (branch_target_d[30]), .\branch_target_d[31] (branch_target_d[31]), 
            .\LM32I_ADR_O[29] (\LM32I_ADR_O[29] ), .\branch_target_d[28] (branch_target_d[28]), 
            .\branch_target_d[29] (branch_target_d[29]), .\LM32I_ADR_O[28] (\LM32I_ADR_O[28] ), 
            .\branch_target_d[26] (branch_target_d[26]), .\branch_target_d[27] (branch_target_d[27]), 
            .\LM32I_ADR_O[27] (\LM32I_ADR_O[27] ), .\branch_target_d[24] (branch_target_d[24]), 
            .\branch_target_d[25] (branch_target_d[25]), .\LM32I_ADR_O[26] (\LM32I_ADR_O[26] ), 
            .\LM32I_ADR_O[25] (\LM32I_ADR_O[25] ), .\branch_target_d[22] (branch_target_d[22]), 
            .\branch_target_d[23] (branch_target_d[23]), .\branch_target_d[20] (branch_target_d[20]), 
            .\branch_target_d[21] (branch_target_d[21]), .\LM32I_ADR_O[24] (\LM32I_ADR_O[24] ), 
            .\LM32I_ADR_O[23] (\LM32I_ADR_O[23] ), .\branch_target_d[18] (branch_target_d[18]), 
            .\branch_target_d[19] (branch_target_d[19]), .\branch_target_d[16] (branch_target_d[16]), 
            .\branch_target_d[17] (branch_target_d[17]), .\LM32I_ADR_O[22] (\LM32I_ADR_O[22] ), 
            .\branch_target_d[14] (branch_target_d[14]), .\branch_target_d[15] (branch_target_d[15]), 
            .\LM32I_ADR_O[21] (\LM32I_ADR_O[21] ), .\branch_target_d[12] (branch_target_d[12]), 
            .\branch_target_d[13] (branch_target_d[13]), .\LM32I_ADR_O[20] (\LM32I_ADR_O[20] ), 
            .\LM32I_ADR_O[19] (\LM32I_ADR_O[19] ), .\LM32I_ADR_O[18] (\LM32I_ADR_O[18] ), 
            .\LM32I_ADR_O[17] (\LM32I_ADR_O[17] ), .\branch_target_d[6] (branch_target_d[6]), 
            .\branch_target_d[7] (branch_target_d[7]), .\LM32I_ADR_O[16] (\LM32I_ADR_O[16] ), 
            .\LM32I_ADR_O[15] (\LM32I_ADR_O[15] ), .\LM32I_ADR_O[14] (\LM32I_ADR_O[14] ), 
            .\branch_target_d[8] (branch_target_d[8]), .\branch_target_d[9] (branch_target_d[9]), 
            .\LM32I_ADR_O[13] (\LM32I_ADR_O[13] ), .\LM32I_ADR_O[12] (\LM32I_ADR_O[12] ), 
            .\branch_target_d[4] (branch_target_d[4]), .\branch_target_d[5] (branch_target_d[5]), 
            .\LM32I_ADR_O[11] (\LM32I_ADR_O[11] ), .\branch_target_d[10] (branch_target_d[10]), 
            .\branch_target_d[11] (branch_target_d[11]), .\LM32I_ADR_O[10] (\LM32I_ADR_O[10] ), 
            .\LM32I_ADR_O[9] (\LM32I_ADR_O[9] ), .\LM32I_ADR_O[8] (\LM32I_ADR_O[8] ), 
            .\LM32I_ADR_O[7] (\LM32I_ADR_O[7] ), .\LM32I_ADR_O[6] (\LM32I_ADR_O[6] ), 
            .\LM32I_ADR_O[5] (\LM32I_ADR_O[5] ), .\LM32I_ADR_O[4] (\LM32I_ADR_O[4] ), 
            .\LM32I_ADR_O[3] (\LM32I_ADR_O[3] ), .n42740(n42740), .n41479(n41479), 
            .n38871(n38871), .w_clk_cpu_enable_878(w_clk_cpu_enable_878), 
            .bus_error_d(bus_error_d), .\instruction_d[31] (instruction_d[31]), 
            .\instruction_d[30] (instruction_d[30]), .\logic_op_d[3] (logic_op_d[3]), 
            .sign_extend_d(instruction[28]), .size_d({size_d}), .read_idx_0_d({read_idx_0_d}), 
            .w_clk_cpu_enable_985(w_clk_cpu_enable_985), .read_idx_1_d({read_idx_1_d}), 
            .\instruction_d[15] (instruction_d[15]), .\instruction_d[14] (instruction_d[14])) /* synthesis syn_module_defined=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(804[5] 896[6])
    \lm32_debug(watchpoints=32'b0)  hw_debug (.dc_re(dc_re), .w_clk_cpu(w_clk_cpu), 
            .dc_re_N_2934(dc_re_N_2934), .\operand_1_x[1] (operand_1_x[1])) /* synthesis syn_module_defined=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1216[5] 1249[6])
    lm32_decoder decoder (.size_d({size_d}), .sign_extend_d(instruction[28]), 
            .\instruction_d[30] (instruction_d[30]), .\instruction_d[31] (instruction_d[31]), 
            .\logic_op_d[3] (logic_op_d[3]), .x_result_sel_csr_d(x_result_sel_csr_d), 
            .\instruction_d[0] (instruction_d[0]), .n1792(n1760[0]), .\instruction_d[15] (instruction_d[15]), 
            .n1777(n1760[15]), .n41397(n41397), .\instruction_d[7] (instruction_d[7]), 
            .n1785(n1760[7]), .\instruction_d[6] (instruction_d[6]), .n1786(n1760[6]), 
            .\instruction_d[5] (instruction_d[5]), .n1787(n1760[5]), .\instruction_d[4] (instruction_d[4]), 
            .n1788(n1760[4]), .\instruction_d[3] (instruction_d[3]), .n1789(n1760[3]), 
            .\instruction_d[2] (instruction_d[2]), .n1790(n1760[2]), .\instruction_d[1] (instruction_d[1]), 
            .n1791(n1760[1]), .n41419(n41419), .n41376(n41376), .adder_op_d_N_1339(adder_op_d_N_1339), 
            .n41361(n41361), .n41364(n41364), .n42740(n42740), .cycles_5__N_2495(cycles_5__N_2495), 
            .n41345(n41345), .n13(n13), .w_clk_cpu_enable_958(w_clk_cpu_enable_958), 
            .n18875(n18875), .x_result_sel_sext_N_1782(x_result_sel_sext_N_1782), 
            .x_bypass_enable_d(x_bypass_enable_d), .m_bypass_enable_d(m_bypass_enable_d), 
            .read_idx_0_d({read_idx_0_d}), .eret_d(eret_d), .bret_d(bret_d), 
            .sign_extend_immediate(sign_extend_immediate), .bus_error_d(bus_error_d), 
            .n41199(n41199), .n41367(n41367), .n41417(n41417), .n22236(n22236), 
            .\instruction_d[12] (instruction_d[12]), .n2(n2_adj_3851), .n2_adj_3(n2_adj_3877), 
            .n2_adj_4(n2_adj_3875), .n2_adj_5(n2_adj_3873), .n2_adj_6(n2_adj_3870), 
            .n2_adj_7(n2_adj_3868), .n2_adj_8(n2_adj_3866), .n2_adj_9(n2_adj_3864), 
            .\instruction_d[8] (instruction_d[8]), .n2_adj_10(n2_adj_3862), 
            .\instruction_d[9] (instruction_d[9]), .n2_adj_11(n2_adj_3858), 
            .\instruction_d[10] (instruction_d[10]), .n2_adj_12(n2_adj_3856), 
            .pc_f({pc_f}), .\bypass_data_0[31] (bypass_data_0[31]), .\d_result_0[31] (d_result_0[31]), 
            .\bypass_data_0[30] (bypass_data_0[30]), .\d_result_0[30] (d_result_0[30]), 
            .\bypass_data_0[29] (bypass_data_0[29]), .\d_result_0[29] (d_result_0[29]), 
            .\bypass_data_0[28] (bypass_data_0[28]), .\d_result_0[28] (d_result_0[28]), 
            .\bypass_data_0[27] (bypass_data_0[27]), .\d_result_0[27] (d_result_0[27]), 
            .n2_adj_13(n2_adj_3879), .\bypass_data_0[26] (bypass_data_0[26]), 
            .\d_result_0[26] (d_result_0[26]), .\bypass_data_0[25] (bypass_data_0[25]), 
            .\d_result_0[25] (d_result_0[25]), .\bypass_data_0[24] (bypass_data_0[24]), 
            .\d_result_0[24] (d_result_0[24]), .\bypass_data_0[23] (bypass_data_0[23]), 
            .\d_result_0[23] (d_result_0[23]), .n22224(n22224), .\instruction_d[11] (instruction_d[11]), 
            .n2_adj_14(n2_adj_3853), .\bypass_data_0[22] (bypass_data_0[22]), 
            .\d_result_0[22] (d_result_0[22]), .\bypass_data_0[21] (bypass_data_0[21]), 
            .\d_result_0[21] (d_result_0[21]), .\bypass_data_0[20] (bypass_data_0[20]), 
            .\d_result_0[20] (d_result_0[20]), .\bypass_data_0[19] (bypass_data_0[19]), 
            .\d_result_0[19] (d_result_0[19]), .\bypass_data_0[18] (bypass_data_0[18]), 
            .\d_result_0[18] (d_result_0[18]), .\bypass_data_0[17] (bypass_data_0[17]), 
            .\d_result_0[17] (d_result_0[17]), .\bypass_data_0[16] (bypass_data_0[16]), 
            .\d_result_0[16] (d_result_0[16]), .\bypass_data_0[15] (bypass_data_0[15]), 
            .\d_result_0[15] (d_result_0[15]), .\bypass_data_0[14] (bypass_data_0[14]), 
            .\d_result_0[14] (d_result_0[14]), .\bypass_data_0[13] (bypass_data_0[13]), 
            .\d_result_0[13] (d_result_0[13]), .\bypass_data_0[12] (bypass_data_0[12]), 
            .\d_result_0[12] (d_result_0[12]), .\bypass_data_0[11] (bypass_data_0[11]), 
            .\d_result_0[11] (d_result_0[11]), .\bypass_data_0[10] (bypass_data_0[10]), 
            .\d_result_0[10] (d_result_0[10]), .\bypass_data_0[9] (bypass_data_0[9]), 
            .\d_result_0[9] (d_result_0[9]), .n42722(n42722), .\bypass_data_0[8] (bypass_data_0[8]), 
            .\d_result_0[8] (d_result_0[8]), .\bypass_data_0[7] (bypass_data_0[7]), 
            .\d_result_0[7] (d_result_0[7]), .\bypass_data_0[6] (bypass_data_0[6]), 
            .\d_result_0[6] (d_result_0[6]), .n41384(n41384), .\bypass_data_0[5] (bypass_data_0[5]), 
            .\d_result_0[5] (d_result_0[5]), .\bypass_data_0[4] (bypass_data_0[4]), 
            .\d_result_0[4] (d_result_0[4]), .n2_adj_15(n2_adj_3842), .\bypass_data_0[3] (bypass_data_0[3]), 
            .\d_result_0[3] (d_result_0[3]), .\instruction_d[14] (instruction_d[14]), 
            .n2_adj_16(n2_adj_3844), .\bypass_data_0[2] (bypass_data_0[2]), 
            .\d_result_0[2] (d_result_0[2]), .\instruction_d[13] (instruction_d[13]), 
            .n2_adj_17(n2_adj_3848), .n41407(n41407), .n1765(n1760[27]), 
            .n1762(n1760[30]), .n1763(n1760[29]), .n1766(n1760[26]), .n1767(n1760[25]), 
            .n1768(n1760[24]), .n1769(n1760[23]), .n1770(n1760[22]), .n1771(n1760[21]), 
            .n1772(n1760[20]), .n1773(n1760[19]), .n1774(n1760[18]), .n1775(n1760[17]), 
            .n1776(n1760[16]), .n1764(n1760[28]), .read_idx_1_d({read_idx_1_d}), 
            .\write_idx_4__N_1770[1] (write_idx_4__N_1770[1]), .bypass_data_1({bypass_data_1}), 
            .n1(n1_adj_3832), .n1_adj_18(n1_adj_3835), .n1_adj_19(n1_adj_3852), 
            .n41394(n41394), .n1_adj_20(n1_adj_3876), .n1_adj_21(n1_adj_3874), 
            .n1_adj_22(n1_adj_3837), .n1_adj_23(n1_adj_3878), .n1_adj_24(n1_adj_3826), 
            .n1_adj_25(n1_adj_3857), .n1_adj_26(n1_adj_3828), .n1_adj_27(n1_adj_3869), 
            .n1_adj_28(n1), .n1_adj_29(n1_adj_3830), .n1_adj_30(n1_adj_3861), 
            .n1_adj_31(n1_adj_3872), .n1_adj_32(n1_adj_3855), .n1_adj_33(n1_adj_3824), 
            .branch_d(branch_d), .n1_adj_34(n1_adj_3882), .n1_adj_35(n1_adj_3867), 
            .n1_adj_36(n1_adj_3886), .n1_adj_37(n1_adj_3850), .n1_adj_38(n1_adj_3839), 
            .n1_adj_39(n1_adj_3820), .n1_adj_40(n1_adj_3843), .n1_adj_41(n1_adj_3863), 
            .n1_adj_42(n1_adj_3847), .n1_adj_43(n1_adj_3888), .n1_adj_44(n1_adj_3841), 
            .n41466(n41466), .x_result_sel_add_N_1785(x_result_sel_add_N_1785), 
            .n1_adj_45(n1_adj_3822), .n1_adj_46(n1_adj_3865), .n1_adj_47(n1_adj_3880), 
            .n1_adj_48(n1_adj_3884), .raw_x_1(raw_x_1), .raw_x_0(raw_x_0), 
            .interlock_N_1327(interlock_N_1327), .n41411(n41411), .raw_m_0(raw_m_0), 
            .interlock_N_1333(interlock_N_1333), .n41406(n41406), .store_d(store_d), 
            .write_enable_N_1809(write_enable_N_1809), .w_result_sel_mul_d(w_result_sel_mul_d), 
            .n25722(n25722), .scall_d(scall_d), .break_d(break_d), .\write_idx_d[4] (write_idx_d[4]), 
            .\write_idx_d[3] (write_idx_d[3]), .\write_idx_d[2] (write_idx_d[2]), 
            .n25724(n25724), .n41380(n41380), .\write_idx_d[0] (write_idx_d[0]), 
            .branch_predict_d(branch_predict_d), .m_result_sel_shift_d(m_result_sel_shift_d)) /* synthesis syn_module_defined=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(899[14] 975[6])
    lm32_adder adder (.muliplicand({muliplicand}), .operand_1_x({operand_1_x}), 
            .adder_op_x(adder_op_x), .adder_op_x_n(adder_op_x_n), .adder_result_x({adder_result_x}), 
            .adder_carry_n_x(adder_carry_n_x)) /* synthesis syn_module_defined=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1046[12] 1056[6])
    
endmodule
//
// Verilog Description of module lm32_shifter
//

module lm32_shifter (left_shift_result, w_clk_cpu, w_clk_cpu_enable_984, 
            \operand_1_x[4] , \operand_1_x[2] , \operand_1_x[3] , direction_m, 
            shifter_result_m, \operand_1_x[1] , \operand_1_x[0] , muliplicand, 
            direction_x, sign_extend_x) /* synthesis syn_module_defined=1 */ ;
    output [31:0]left_shift_result;
    input w_clk_cpu;
    input w_clk_cpu_enable_984;
    input \operand_1_x[4] ;
    input \operand_1_x[2] ;
    input \operand_1_x[3] ;
    output direction_m;
    output [31:0]shifter_result_m;
    input \operand_1_x[1] ;
    input \operand_1_x[0] ;
    input [31:0]muliplicand;
    input direction_x;
    input sign_extend_x;
    
    wire w_clk_cpu /* synthesis SET_AS_NETWORK=w_clk_cpu, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(22[6:15])
    wire [63:0]left_shift_result_31__N_2188;
    
    wire n41339, n211, n41337, n71, n41338, n41333, n212, n41331, 
        n72, n41332, n41328, n141, n41329, n41325, n143, n41326, 
        n41322, n144, n41323, n41287, n138, n41288, n41285, n4, 
        n41286, n41798, n3, n41799, n41282, n142, n41283, n39751, 
        n39752, n39754, n39755, n39757, n39758, n208, n224, n207, 
        n223;
    wire [31:0]right_shift_operand;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(96[23:42])
    
    wire n206, n222, n205, n221, n70, n41441, fill_value, n210, 
        n41801, n209, n69, n41800, n41797, n41414, n31, n41440, 
        n154, n39779, n146, n39778, n6, n8, n10, n12, n74, 
        n150, n158, n214, n156, n94, n155, n153, n78, n82, 
        n86, n90, n5, n7, n216, n152, n160, n215, n151, n159, 
        n213, n149, n157, n93, n148, n147, n145, n9, n137, 
        n73, n77, n81, n85, n17, n19, n21, n23, n11, n13, 
        n15, n89, n25, n27, n29, n75, n79, n139, n83, n87, 
        n91, n95, n76, n80, n140, n84, n88, n20, n22, n24, 
        n26, n14, n16, n18, n92, n96, n28, n30, n32, n41481, 
        n41482, n41480;
    
    FD1P3AX right_shift_result_i0_i11 (.D(left_shift_result_31__N_2188[11]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[20])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i11.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i10 (.D(left_shift_result_31__N_2188[10]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[21])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i10.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i9 (.D(left_shift_result_31__N_2188[9]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[22])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i9.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i8 (.D(left_shift_result_31__N_2188[8]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[23])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i8.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i7 (.D(left_shift_result_31__N_2188[7]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[24])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i7.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i6 (.D(left_shift_result_31__N_2188[6]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[25])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i6.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i5 (.D(left_shift_result_31__N_2188[5]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[26])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i5.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i4 (.D(left_shift_result_31__N_2188[4]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[27])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i4.GSR = "ENABLED";
    PFUMX i38563 (.BLUT(n41339), .ALUT(n211), .C0(\operand_1_x[4] ), .Z(left_shift_result_31__N_2188[2]));
    FD1P3AX right_shift_result_i0_i3 (.D(left_shift_result_31__N_2188[3]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[28])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i3.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i2 (.D(left_shift_result_31__N_2188[2]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[29])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i2.GSR = "ENABLED";
    PFUMX i38561 (.BLUT(n41337), .ALUT(n71), .C0(\operand_1_x[2] ), .Z(n41338));
    FD1P3AX right_shift_result_i0_i1 (.D(left_shift_result_31__N_2188[1]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[30])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i1.GSR = "ENABLED";
    PFUMX i38559 (.BLUT(n41333), .ALUT(n212), .C0(\operand_1_x[4] ), .Z(left_shift_result_31__N_2188[3]));
    PFUMX i38557 (.BLUT(n41331), .ALUT(n72), .C0(\operand_1_x[2] ), .Z(n41332));
    PFUMX i38555 (.BLUT(n41328), .ALUT(n141), .C0(\operand_1_x[3] ), .Z(n41329));
    PFUMX i38553 (.BLUT(n41325), .ALUT(n143), .C0(\operand_1_x[3] ), .Z(n41326));
    PFUMX i38551 (.BLUT(n41322), .ALUT(n144), .C0(\operand_1_x[3] ), .Z(n41323));
    LUT4 left_shift_result_0__I_0_21_i2_3_lut (.A(left_shift_result[30]), 
         .B(left_shift_result[1]), .C(direction_m), .Z(shifter_result_m[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i2_3_lut.init = 16'hcaca;
    FD1P3AX right_shift_result_i0_i0 (.D(left_shift_result_31__N_2188[0]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[31])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i0.GSR = "ENABLED";
    PFUMX i38520 (.BLUT(n41287), .ALUT(n138), .C0(\operand_1_x[3] ), .Z(n41288));
    PFUMX i38518 (.BLUT(n41285), .ALUT(n4), .C0(\operand_1_x[1] ), .Z(n41286));
    LUT4 n41798_bdd_3_lut (.A(n41798), .B(n3), .C(\operand_1_x[1] ), .Z(n41799)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41798_bdd_3_lut.init = 16'hcaca;
    PFUMX i38516 (.BLUT(n41282), .ALUT(n142), .C0(\operand_1_x[3] ), .Z(n41283));
    PFUMX i37199 (.BLUT(n39751), .ALUT(n39752), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2188[8]));
    PFUMX i37202 (.BLUT(n39754), .ALUT(n39755), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2188[10]));
    PFUMX i37205 (.BLUT(n39757), .ALUT(n39758), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2188[11]));
    PFUMX shift_right_13_i272 (.BLUT(n208), .ALUT(n224), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2188[15])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;
    PFUMX shift_right_13_i271 (.BLUT(n207), .ALUT(n223), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2188[14])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;
    LUT4 n4_bdd_3_lut_38768 (.A(right_shift_operand[2]), .B(right_shift_operand[1]), 
         .C(\operand_1_x[0] ), .Z(n41285)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n4_bdd_3_lut_38768.init = 16'hacac;
    PFUMX shift_right_13_i270 (.BLUT(n206), .ALUT(n222), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2188[13])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;
    PFUMX shift_right_13_i269 (.BLUT(n205), .ALUT(n221), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2188[12])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;
    LUT4 n41286_bdd_3_lut (.A(n41286), .B(n70), .C(\operand_1_x[2] ), 
         .Z(n41287)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41286_bdd_3_lut.init = 16'hcaca;
    LUT4 i21448_3_lut_4_lut (.A(n41441), .B(\operand_1_x[3] ), .C(fill_value), 
         .D(right_shift_operand[31]), .Z(n224)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i21448_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n41288_bdd_3_lut (.A(n41288), .B(n210), .C(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2188[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41288_bdd_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i3_3_lut (.A(left_shift_result[29]), 
         .B(left_shift_result[2]), .C(direction_m), .Z(shifter_result_m[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i3_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i4_3_lut (.A(left_shift_result[28]), 
         .B(left_shift_result[3]), .C(direction_m), .Z(shifter_result_m[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i4_3_lut.init = 16'hcaca;
    PFUMX i38733 (.BLUT(n41801), .ALUT(n209), .C0(\operand_1_x[4] ), .Z(left_shift_result_31__N_2188[0]));
    PFUMX i38731 (.BLUT(n41799), .ALUT(n69), .C0(\operand_1_x[2] ), .Z(n41800));
    PFUMX i38729 (.BLUT(n41797), .ALUT(right_shift_operand[1]), .C0(\operand_1_x[0] ), 
          .Z(n41798));
    LUT4 left_shift_result_0__I_0_21_i1_3_lut (.A(left_shift_result[31]), 
         .B(left_shift_result[0]), .C(direction_m), .Z(shifter_result_m[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i1_3_lut.init = 16'hcaca;
    LUT4 i21466_4_lut (.A(right_shift_operand[31]), .B(fill_value), .C(n41414), 
         .D(\operand_1_x[4] ), .Z(left_shift_result_31__N_2188[31])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i21466_4_lut.init = 16'hccca;
    LUT4 i21464_4_lut (.A(n31), .B(fill_value), .C(n41440), .D(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2188[30])) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i21464_4_lut.init = 16'hccca;
    LUT4 i37225_3_lut (.A(n154), .B(fill_value), .C(\operand_1_x[3] ), 
         .Z(n39779)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37225_3_lut.init = 16'hcaca;
    LUT4 i37224_3_lut (.A(n138), .B(n146), .C(\operand_1_x[3] ), .Z(n39778)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37224_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i70_3_lut (.A(n6), .B(n8), .C(\operand_1_x[1] ), 
         .Z(n70)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i70_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i74_3_lut (.A(n10), .B(n12), .C(\operand_1_x[1] ), 
         .Z(n74)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i74_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i10_3_lut (.A(right_shift_operand[9]), .B(right_shift_operand[10]), 
         .C(\operand_1_x[0] ), .Z(n10)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i10_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i6_3_lut (.A(right_shift_operand[5]), .B(right_shift_operand[6]), 
         .C(\operand_1_x[0] ), .Z(n6)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i6_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i8_3_lut (.A(right_shift_operand[7]), .B(right_shift_operand[8]), 
         .C(\operand_1_x[0] ), .Z(n8)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i8_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i8_3_lut (.A(muliplicand[7]), .B(muliplicand[24]), 
         .C(direction_x), .Z(right_shift_operand[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i8_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i6_3_lut (.A(muliplicand[5]), .B(muliplicand[26]), 
         .C(direction_x), .Z(right_shift_operand[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i6_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i7_3_lut (.A(muliplicand[6]), .B(muliplicand[25]), 
         .C(direction_x), .Z(right_shift_operand[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i7_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i214_3_lut (.A(n150), .B(n158), .C(\operand_1_x[3] ), 
         .Z(n214)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i214_3_lut.init = 16'hcaca;
    LUT4 i21458_3_lut_4_lut (.A(\operand_1_x[3] ), .B(\operand_1_x[4] ), 
         .C(fill_value), .D(n156), .Z(left_shift_result_31__N_2188[27])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i21458_3_lut_4_lut.init = 16'hf1e0;
    LUT4 shift_right_13_i158_3_lut (.A(n94), .B(fill_value), .C(\operand_1_x[2] ), 
         .Z(n158)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i158_3_lut.init = 16'hcaca;
    LUT4 i21454_3_lut_4_lut (.A(\operand_1_x[3] ), .B(\operand_1_x[4] ), 
         .C(fill_value), .D(n154), .Z(left_shift_result_31__N_2188[25])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i21454_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i21456_3_lut_4_lut (.A(\operand_1_x[3] ), .B(\operand_1_x[4] ), 
         .C(fill_value), .D(n155), .Z(left_shift_result_31__N_2188[26])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i21456_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i21452_3_lut_4_lut (.A(\operand_1_x[3] ), .B(\operand_1_x[4] ), 
         .C(fill_value), .D(n153), .Z(left_shift_result_31__N_2188[24])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i21452_3_lut_4_lut.init = 16'hf1e0;
    LUT4 shift_right_13_i138_3_lut (.A(n74), .B(n78), .C(\operand_1_x[2] ), 
         .Z(n138)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i138_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i4_3_lut (.A(right_shift_operand[3]), .B(right_shift_operand[4]), 
         .C(\operand_1_x[0] ), .Z(n4)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i4_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i4_3_lut (.A(muliplicand[3]), .B(muliplicand[28]), 
         .C(direction_x), .Z(right_shift_operand[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i4_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i5_3_lut (.A(muliplicand[4]), .B(muliplicand[27]), 
         .C(direction_x), .Z(right_shift_operand[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i5_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i210_3_lut (.A(n146), .B(n154), .C(\operand_1_x[3] ), 
         .Z(n210)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i210_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i146_3_lut (.A(n82), .B(n86), .C(\operand_1_x[2] ), 
         .Z(n146)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i146_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i154_3_lut (.A(n90), .B(n94), .C(\operand_1_x[2] ), 
         .Z(n154)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i154_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i2_3_lut (.A(muliplicand[1]), .B(muliplicand[30]), 
         .C(direction_x), .Z(right_shift_operand[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i2_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i3_3_lut (.A(muliplicand[2]), .B(muliplicand[29]), 
         .C(direction_x), .Z(right_shift_operand[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i3_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i5_3_lut (.A(left_shift_result[27]), 
         .B(left_shift_result[4]), .C(direction_m), .Z(shifter_result_m[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i5_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i69_3_lut (.A(n5), .B(n7), .C(\operand_1_x[1] ), 
         .Z(n69)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i69_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i5_3_lut (.A(right_shift_operand[4]), .B(right_shift_operand[5]), 
         .C(\operand_1_x[0] ), .Z(n5)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i5_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i7_3_lut (.A(right_shift_operand[6]), .B(right_shift_operand[7]), 
         .C(\operand_1_x[0] ), .Z(n7)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i7_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i3_3_lut (.A(right_shift_operand[2]), .B(right_shift_operand[3]), 
         .C(\operand_1_x[0] ), .Z(n3)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i3_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i280_3_lut (.A(n216), .B(fill_value), .C(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2188[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i280_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i216_3_lut (.A(n152), .B(n160), .C(\operand_1_x[3] ), 
         .Z(n216)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i216_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i279_3_lut (.A(n215), .B(fill_value), .C(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2188[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i279_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i215_3_lut (.A(n151), .B(n159), .C(\operand_1_x[3] ), 
         .Z(n215)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i215_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i278_3_lut (.A(n214), .B(fill_value), .C(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2188[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i278_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i6_3_lut (.A(left_shift_result[26]), 
         .B(left_shift_result[5]), .C(direction_m), .Z(shifter_result_m[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i6_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i277_3_lut (.A(n213), .B(fill_value), .C(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2188[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i277_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i213_3_lut (.A(n149), .B(n157), .C(\operand_1_x[3] ), 
         .Z(n213)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i213_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i157_3_lut (.A(n93), .B(fill_value), .C(\operand_1_x[2] ), 
         .Z(n157)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i157_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i276_3_lut (.A(n212), .B(fill_value), .C(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2188[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i276_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i212_3_lut (.A(n148), .B(n156), .C(\operand_1_x[3] ), 
         .Z(n212)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i212_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i275_3_lut (.A(n211), .B(fill_value), .C(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2188[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i275_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i211_3_lut (.A(n147), .B(n155), .C(\operand_1_x[3] ), 
         .Z(n211)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i211_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i274_3_lut (.A(n210), .B(fill_value), .C(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2188[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i274_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i273_3_lut (.A(n209), .B(fill_value), .C(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2188[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i273_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i209_3_lut (.A(n145), .B(n153), .C(\operand_1_x[3] ), 
         .Z(n209)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i209_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i72_3_lut (.A(n8), .B(n10), .C(\operand_1_x[1] ), 
         .Z(n72)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i72_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i71_3_lut (.A(n7), .B(n9), .C(\operand_1_x[1] ), 
         .Z(n71)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i71_3_lut.init = 16'hcaca;
    LUT4 right_shift_operand_1__bdd_3_lut_38735 (.A(muliplicand[31]), .B(muliplicand[0]), 
         .C(direction_x), .Z(n41797)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam right_shift_operand_1__bdd_3_lut_38735.init = 16'hacac;
    LUT4 n41800_bdd_3_lut (.A(n41800), .B(n137), .C(\operand_1_x[3] ), 
         .Z(n41801)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41800_bdd_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i137_3_lut (.A(n73), .B(n77), .C(\operand_1_x[2] ), 
         .Z(n137)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i137_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i145_3_lut (.A(n81), .B(n85), .C(\operand_1_x[2] ), 
         .Z(n145)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i145_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i81_3_lut (.A(n17), .B(n19), .C(\operand_1_x[1] ), 
         .Z(n81)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i81_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i85_3_lut (.A(n21), .B(n23), .C(\operand_1_x[1] ), 
         .Z(n85)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i85_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i21_3_lut (.A(right_shift_operand[20]), .B(right_shift_operand[21]), 
         .C(\operand_1_x[0] ), .Z(n21)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i21_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i23_3_lut (.A(right_shift_operand[22]), .B(right_shift_operand[23]), 
         .C(\operand_1_x[0] ), .Z(n23)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i23_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i23_3_lut (.A(muliplicand[22]), .B(muliplicand[9]), 
         .C(direction_x), .Z(right_shift_operand[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i23_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i24_3_lut (.A(muliplicand[23]), .B(muliplicand[8]), 
         .C(direction_x), .Z(right_shift_operand[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i24_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i21_3_lut (.A(muliplicand[20]), .B(muliplicand[11]), 
         .C(direction_x), .Z(right_shift_operand[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i21_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i22_3_lut (.A(muliplicand[21]), .B(muliplicand[10]), 
         .C(direction_x), .Z(right_shift_operand[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i22_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i73_3_lut (.A(n9), .B(n11), .C(\operand_1_x[1] ), 
         .Z(n73)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i73_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i77_3_lut (.A(n13), .B(n15), .C(\operand_1_x[1] ), 
         .Z(n77)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i77_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i13_3_lut (.A(right_shift_operand[12]), .B(right_shift_operand[13]), 
         .C(\operand_1_x[0] ), .Z(n13)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i13_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i15_3_lut (.A(right_shift_operand[14]), .B(right_shift_operand[15]), 
         .C(\operand_1_x[0] ), .Z(n15)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i15_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i16_3_lut (.A(muliplicand[15]), .B(muliplicand[16]), 
         .C(direction_x), .Z(right_shift_operand[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i16_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i9_3_lut (.A(right_shift_operand[8]), .B(right_shift_operand[9]), 
         .C(\operand_1_x[0] ), .Z(n9)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i9_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i11_3_lut (.A(right_shift_operand[10]), .B(right_shift_operand[11]), 
         .C(\operand_1_x[0] ), .Z(n11)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i11_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i9_3_lut (.A(muliplicand[8]), .B(muliplicand[23]), 
         .C(direction_x), .Z(right_shift_operand[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i9_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i10_3_lut (.A(muliplicand[9]), .B(muliplicand[22]), 
         .C(direction_x), .Z(right_shift_operand[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i10_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i11_3_lut (.A(muliplicand[10]), .B(muliplicand[21]), 
         .C(direction_x), .Z(right_shift_operand[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i11_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i12_3_lut (.A(muliplicand[11]), .B(muliplicand[20]), 
         .C(direction_x), .Z(right_shift_operand[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i12_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i15_3_lut (.A(muliplicand[14]), .B(muliplicand[17]), 
         .C(direction_x), .Z(right_shift_operand[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i15_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i13_3_lut (.A(muliplicand[12]), .B(muliplicand[19]), 
         .C(direction_x), .Z(right_shift_operand[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i13_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i14_3_lut (.A(muliplicand[13]), .B(muliplicand[18]), 
         .C(direction_x), .Z(right_shift_operand[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i14_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i17_3_lut (.A(right_shift_operand[16]), .B(right_shift_operand[17]), 
         .C(\operand_1_x[0] ), .Z(n17)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i17_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i17_3_lut (.A(muliplicand[16]), .B(muliplicand[15]), 
         .C(direction_x), .Z(right_shift_operand[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i17_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i19_3_lut (.A(right_shift_operand[18]), .B(right_shift_operand[19]), 
         .C(\operand_1_x[0] ), .Z(n19)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i19_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i18_3_lut (.A(muliplicand[17]), .B(muliplicand[14]), 
         .C(direction_x), .Z(right_shift_operand[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i18_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i19_3_lut (.A(muliplicand[18]), .B(muliplicand[13]), 
         .C(direction_x), .Z(right_shift_operand[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i19_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i20_3_lut (.A(muliplicand[19]), .B(muliplicand[12]), 
         .C(direction_x), .Z(right_shift_operand[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i20_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i153_3_lut (.A(n89), .B(n93), .C(\operand_1_x[2] ), 
         .Z(n153)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i153_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut (.A(direction_x), .B(muliplicand[31]), .C(sign_extend_x), 
         .Z(fill_value)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(116[21] 118[29])
    defparam i2_3_lut.init = 16'h4040;
    LUT4 shift_right_13_i89_3_lut (.A(n25), .B(n27), .C(\operand_1_x[1] ), 
         .Z(n89)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i89_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i93_3_lut (.A(n29), .B(n31), .C(\operand_1_x[1] ), 
         .Z(n93)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i93_3_lut.init = 16'hcaca;
    LUT4 n142_bdd_3_lut (.A(n70), .B(n74), .C(\operand_1_x[2] ), .Z(n41282)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n142_bdd_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i25_3_lut (.A(right_shift_operand[24]), .B(right_shift_operand[25]), 
         .C(\operand_1_x[0] ), .Z(n25)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i25_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i27_3_lut (.A(right_shift_operand[26]), .B(right_shift_operand[27]), 
         .C(\operand_1_x[0] ), .Z(n27)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i27_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i25_3_lut (.A(muliplicand[24]), .B(muliplicand[7]), 
         .C(direction_x), .Z(right_shift_operand[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i25_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i26_3_lut (.A(muliplicand[25]), .B(muliplicand[6]), 
         .C(direction_x), .Z(right_shift_operand[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i26_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i27_3_lut (.A(muliplicand[26]), .B(muliplicand[5]), 
         .C(direction_x), .Z(right_shift_operand[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i27_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i28_3_lut (.A(muliplicand[27]), .B(muliplicand[4]), 
         .C(direction_x), .Z(right_shift_operand[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i28_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i29_3_lut (.A(right_shift_operand[28]), .B(right_shift_operand[29]), 
         .C(\operand_1_x[0] ), .Z(n29)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i29_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i31_3_lut (.A(right_shift_operand[30]), .B(right_shift_operand[31]), 
         .C(\operand_1_x[0] ), .Z(n31)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i31_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i31_3_lut (.A(muliplicand[30]), .B(muliplicand[1]), 
         .C(direction_x), .Z(right_shift_operand[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i31_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i32_3_lut (.A(muliplicand[31]), .B(muliplicand[0]), 
         .C(direction_x), .Z(right_shift_operand[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i32_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i29_3_lut (.A(muliplicand[28]), .B(muliplicand[3]), 
         .C(direction_x), .Z(right_shift_operand[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i29_3_lut.init = 16'hcaca;
    LUT4 operand_0_x_31__I_0_22_i30_3_lut (.A(muliplicand[29]), .B(muliplicand[2]), 
         .C(direction_x), .Z(right_shift_operand[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(113[30:99])
    defparam operand_0_x_31__I_0_22_i30_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i139_3_lut (.A(n75), .B(n79), .C(\operand_1_x[2] ), 
         .Z(n139)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i139_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i147_3_lut (.A(n83), .B(n87), .C(\operand_1_x[2] ), 
         .Z(n147)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i147_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i83_3_lut (.A(n19), .B(n21), .C(\operand_1_x[1] ), 
         .Z(n83)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i83_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i87_3_lut (.A(n23), .B(n25), .C(\operand_1_x[1] ), 
         .Z(n87)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i87_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i75_3_lut (.A(n11), .B(n13), .C(\operand_1_x[1] ), 
         .Z(n75)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i75_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i79_3_lut (.A(n15), .B(n17), .C(\operand_1_x[1] ), 
         .Z(n79)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i79_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i155_3_lut (.A(n91), .B(n95), .C(\operand_1_x[2] ), 
         .Z(n155)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i155_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i95_3_lut (.A(n31), .B(fill_value), .C(\operand_1_x[1] ), 
         .Z(n95)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i95_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i91_3_lut (.A(n27), .B(n29), .C(\operand_1_x[1] ), 
         .Z(n91)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i91_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i140_3_lut (.A(n76), .B(n80), .C(\operand_1_x[2] ), 
         .Z(n140)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i140_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i148_3_lut (.A(n84), .B(n88), .C(\operand_1_x[2] ), 
         .Z(n148)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i148_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i84_3_lut (.A(n20), .B(n22), .C(\operand_1_x[1] ), 
         .Z(n84)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i84_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i88_3_lut (.A(n24), .B(n26), .C(\operand_1_x[1] ), 
         .Z(n88)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i88_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i24_3_lut (.A(right_shift_operand[23]), .B(right_shift_operand[24]), 
         .C(\operand_1_x[0] ), .Z(n24)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i24_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i26_3_lut (.A(right_shift_operand[25]), .B(right_shift_operand[26]), 
         .C(\operand_1_x[0] ), .Z(n26)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i26_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i76_3_lut (.A(n12), .B(n14), .C(\operand_1_x[1] ), 
         .Z(n76)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i76_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i80_3_lut (.A(n16), .B(n18), .C(\operand_1_x[1] ), 
         .Z(n80)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i80_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i16_4_lut (.A(muliplicand[15]), .B(muliplicand[16]), 
         .C(direction_x), .D(\operand_1_x[0] ), .Z(n16)) /* synthesis lut_function=(A (B+(C (D)+!C !(D)))+!A !((C (D)+!C !(D))+!B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i16_4_lut.init = 16'hacca;
    LUT4 shift_right_13_i18_3_lut (.A(right_shift_operand[17]), .B(right_shift_operand[18]), 
         .C(\operand_1_x[0] ), .Z(n18)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i18_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i12_3_lut (.A(right_shift_operand[11]), .B(right_shift_operand[12]), 
         .C(\operand_1_x[0] ), .Z(n12)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i12_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i14_3_lut (.A(right_shift_operand[13]), .B(right_shift_operand[14]), 
         .C(\operand_1_x[0] ), .Z(n14)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i14_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i20_3_lut (.A(right_shift_operand[19]), .B(right_shift_operand[20]), 
         .C(\operand_1_x[0] ), .Z(n20)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i20_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i22_3_lut (.A(right_shift_operand[21]), .B(right_shift_operand[22]), 
         .C(\operand_1_x[0] ), .Z(n22)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i22_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i156_3_lut (.A(n92), .B(n96), .C(\operand_1_x[2] ), 
         .Z(n156)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i156_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i92_3_lut (.A(n28), .B(n30), .C(\operand_1_x[1] ), 
         .Z(n92)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i92_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i28_3_lut (.A(right_shift_operand[27]), .B(right_shift_operand[28]), 
         .C(\operand_1_x[0] ), .Z(n28)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i28_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i30_3_lut (.A(right_shift_operand[29]), .B(right_shift_operand[30]), 
         .C(\operand_1_x[0] ), .Z(n30)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i30_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i144_3_lut (.A(n80), .B(n84), .C(\operand_1_x[2] ), 
         .Z(n144)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i144_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i152_3_lut (.A(n88), .B(n92), .C(\operand_1_x[2] ), 
         .Z(n152)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i152_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i143_3_lut (.A(n79), .B(n83), .C(\operand_1_x[2] ), 
         .Z(n143)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i143_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i151_3_lut (.A(n87), .B(n91), .C(\operand_1_x[2] ), 
         .Z(n151)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i151_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i142_3_lut (.A(n78), .B(n82), .C(\operand_1_x[2] ), 
         .Z(n142)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i142_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i150_3_lut (.A(n86), .B(n90), .C(\operand_1_x[2] ), 
         .Z(n150)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i150_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i86_3_lut (.A(n22), .B(n24), .C(\operand_1_x[1] ), 
         .Z(n86)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i86_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i90_3_lut (.A(n26), .B(n28), .C(\operand_1_x[1] ), 
         .Z(n90)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i90_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i78_3_lut (.A(n14), .B(n16), .C(\operand_1_x[1] ), 
         .Z(n78)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i78_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i82_3_lut (.A(n18), .B(n20), .C(\operand_1_x[1] ), 
         .Z(n82)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i82_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i94_3_lut (.A(n30), .B(n32), .C(\operand_1_x[1] ), 
         .Z(n94)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i94_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i32_3_lut (.A(right_shift_operand[31]), .B(fill_value), 
         .C(\operand_1_x[0] ), .Z(n32)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i32_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i141_3_lut (.A(n77), .B(n81), .C(\operand_1_x[2] ), 
         .Z(n141)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i141_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i149_3_lut (.A(n85), .B(n89), .C(\operand_1_x[2] ), 
         .Z(n149)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i149_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i205_3_lut (.A(n141), .B(n149), .C(\operand_1_x[3] ), 
         .Z(n205)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i205_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i206_3_lut (.A(n142), .B(n150), .C(\operand_1_x[3] ), 
         .Z(n206)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i206_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i207_3_lut (.A(n143), .B(n151), .C(\operand_1_x[3] ), 
         .Z(n207)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i207_3_lut.init = 16'hcaca;
    LUT4 shift_right_13_i208_3_lut (.A(n144), .B(n152), .C(\operand_1_x[3] ), 
         .Z(n208)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam shift_right_13_i208_3_lut.init = 16'hcaca;
    LUT4 i37204_3_lut (.A(n156), .B(fill_value), .C(\operand_1_x[3] ), 
         .Z(n39758)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37204_3_lut.init = 16'hcaca;
    LUT4 i37203_3_lut (.A(n140), .B(n148), .C(\operand_1_x[3] ), .Z(n39757)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37203_3_lut.init = 16'hcaca;
    LUT4 i37201_3_lut (.A(n155), .B(fill_value), .C(\operand_1_x[3] ), 
         .Z(n39755)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37201_3_lut.init = 16'hcaca;
    LUT4 i37200_3_lut (.A(n139), .B(n147), .C(\operand_1_x[3] ), .Z(n39754)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37200_3_lut.init = 16'hcaca;
    LUT4 i21446_3_lut_4_lut (.A(n41481), .B(\operand_1_x[3] ), .C(fill_value), 
         .D(n31), .Z(n223)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i21446_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i37198_3_lut (.A(n153), .B(fill_value), .C(\operand_1_x[3] ), 
         .Z(n39752)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37198_3_lut.init = 16'hcaca;
    LUT4 i37197_3_lut (.A(n137), .B(n145), .C(\operand_1_x[3] ), .Z(n39751)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37197_3_lut.init = 16'hcaca;
    LUT4 i21423_3_lut_4_lut (.A(n41482), .B(\operand_1_x[2] ), .C(fill_value), 
         .D(right_shift_operand[31]), .Z(n160)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i21423_3_lut_4_lut.init = 16'hf1e0;
    LUT4 n41283_bdd_3_lut (.A(n41283), .B(n214), .C(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2188[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41283_bdd_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i7_3_lut (.A(left_shift_result[25]), 
         .B(left_shift_result[6]), .C(direction_m), .Z(shifter_result_m[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i7_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i8_3_lut (.A(left_shift_result[24]), 
         .B(left_shift_result[7]), .C(direction_m), .Z(shifter_result_m[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i8_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i9_3_lut (.A(left_shift_result[23]), 
         .B(left_shift_result[8]), .C(direction_m), .Z(shifter_result_m[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i9_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i10_3_lut (.A(left_shift_result[22]), 
         .B(left_shift_result[9]), .C(direction_m), .Z(shifter_result_m[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i10_3_lut.init = 16'hcaca;
    LUT4 i21462_3_lut_4_lut (.A(n41480), .B(\operand_1_x[4] ), .C(fill_value), 
         .D(n94), .Z(left_shift_result_31__N_2188[29])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i21462_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i21460_3_lut_4_lut (.A(n41480), .B(\operand_1_x[4] ), .C(fill_value), 
         .D(n93), .Z(left_shift_result_31__N_2188[28])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i21460_3_lut_4_lut.init = 16'hf1e0;
    LUT4 left_shift_result_0__I_0_21_i11_3_lut (.A(left_shift_result[21]), 
         .B(left_shift_result[10]), .C(direction_m), .Z(shifter_result_m[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i11_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i12_3_lut (.A(left_shift_result[20]), 
         .B(left_shift_result[11]), .C(direction_m), .Z(shifter_result_m[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i12_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i13_3_lut (.A(left_shift_result[19]), 
         .B(left_shift_result[12]), .C(direction_m), .Z(shifter_result_m[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i13_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i14_3_lut (.A(left_shift_result[18]), 
         .B(left_shift_result[13]), .C(direction_m), .Z(shifter_result_m[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i14_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i15_3_lut (.A(left_shift_result[17]), 
         .B(left_shift_result[14]), .C(direction_m), .Z(shifter_result_m[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i15_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i16_3_lut (.A(left_shift_result[16]), 
         .B(left_shift_result[15]), .C(direction_m), .Z(shifter_result_m[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i16_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i17_3_lut (.A(left_shift_result[15]), 
         .B(left_shift_result[16]), .C(direction_m), .Z(shifter_result_m[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i17_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i18_3_lut (.A(left_shift_result[14]), 
         .B(left_shift_result[17]), .C(direction_m), .Z(shifter_result_m[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i18_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i19_3_lut (.A(left_shift_result[13]), 
         .B(left_shift_result[18]), .C(direction_m), .Z(shifter_result_m[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i19_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i20_3_lut (.A(left_shift_result[12]), 
         .B(left_shift_result[19]), .C(direction_m), .Z(shifter_result_m[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i20_3_lut.init = 16'hcaca;
    FD1P3AX direction_m_20 (.D(direction_x), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(direction_m));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam direction_m_20.GSR = "ENABLED";
    LUT4 left_shift_result_0__I_0_21_i21_3_lut (.A(left_shift_result[11]), 
         .B(left_shift_result[20]), .C(direction_m), .Z(shifter_result_m[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i21_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i22_3_lut (.A(left_shift_result[10]), 
         .B(left_shift_result[21]), .C(direction_m), .Z(shifter_result_m[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i22_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i23_3_lut (.A(left_shift_result[9]), 
         .B(left_shift_result[22]), .C(direction_m), .Z(shifter_result_m[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i23_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i24_3_lut (.A(left_shift_result[8]), 
         .B(left_shift_result[23]), .C(direction_m), .Z(shifter_result_m[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i24_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i25_3_lut (.A(left_shift_result[7]), 
         .B(left_shift_result[24]), .C(direction_m), .Z(shifter_result_m[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i25_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i26_3_lut (.A(left_shift_result[6]), 
         .B(left_shift_result[25]), .C(direction_m), .Z(shifter_result_m[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i26_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i27_3_lut (.A(left_shift_result[5]), 
         .B(left_shift_result[26]), .C(direction_m), .Z(shifter_result_m[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i27_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i28_3_lut (.A(left_shift_result[4]), 
         .B(left_shift_result[27]), .C(direction_m), .Z(shifter_result_m[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i28_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i29_3_lut (.A(left_shift_result[3]), 
         .B(left_shift_result[28]), .C(direction_m), .Z(shifter_result_m[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i29_3_lut.init = 16'hcaca;
    LUT4 n144_bdd_3_lut_38791 (.A(n72), .B(n76), .C(\operand_1_x[2] ), 
         .Z(n41322)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n144_bdd_3_lut_38791.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i30_3_lut (.A(left_shift_result[2]), 
         .B(left_shift_result[29]), .C(direction_m), .Z(shifter_result_m[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i30_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i31_3_lut (.A(left_shift_result[1]), 
         .B(left_shift_result[30]), .C(direction_m), .Z(shifter_result_m[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i31_3_lut.init = 16'hcaca;
    LUT4 left_shift_result_0__I_0_21_i32_3_lut (.A(left_shift_result[0]), 
         .B(left_shift_result[31]), .C(direction_m), .Z(shifter_result_m[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(131[27:102])
    defparam left_shift_result_0__I_0_21_i32_3_lut.init = 16'hcaca;
    LUT4 n41323_bdd_3_lut (.A(n41323), .B(n216), .C(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2188[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41323_bdd_3_lut.init = 16'hcaca;
    LUT4 n143_bdd_3_lut_38794 (.A(n71), .B(n75), .C(\operand_1_x[2] ), 
         .Z(n41325)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n143_bdd_3_lut_38794.init = 16'hcaca;
    LUT4 n41326_bdd_3_lut (.A(n41326), .B(n215), .C(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2188[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41326_bdd_3_lut.init = 16'hcaca;
    LUT4 n141_bdd_3_lut (.A(n69), .B(n73), .C(\operand_1_x[2] ), .Z(n41328)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n141_bdd_3_lut.init = 16'hcaca;
    LUT4 n41329_bdd_3_lut (.A(n41329), .B(n213), .C(\operand_1_x[4] ), 
         .Z(left_shift_result_31__N_2188[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41329_bdd_3_lut.init = 16'hcaca;
    LUT4 n72_bdd_3_lut (.A(n4), .B(n6), .C(\operand_1_x[1] ), .Z(n41331)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n72_bdd_3_lut.init = 16'hcaca;
    LUT4 n41332_bdd_3_lut (.A(n41332), .B(n140), .C(\operand_1_x[3] ), 
         .Z(n41333)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41332_bdd_3_lut.init = 16'hcaca;
    FD1P3AX right_shift_result_i0_i31 (.D(left_shift_result_31__N_2188[31]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i31.GSR = "ENABLED";
    LUT4 n71_bdd_3_lut (.A(n3), .B(n5), .C(\operand_1_x[1] ), .Z(n41337)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n71_bdd_3_lut.init = 16'hcaca;
    LUT4 n41338_bdd_3_lut (.A(n41338), .B(n139), .C(\operand_1_x[3] ), 
         .Z(n41339)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41338_bdd_3_lut.init = 16'hcaca;
    FD1P3AX right_shift_result_i0_i30 (.D(left_shift_result_31__N_2188[30]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i30.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i29 (.D(left_shift_result_31__N_2188[29]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i29.GSR = "ENABLED";
    LUT4 i21441_2_lut_rep_393 (.A(\operand_1_x[2] ), .B(\operand_1_x[3] ), 
         .Z(n41480)) /* synthesis lut_function=(A+(B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i21441_2_lut_rep_393.init = 16'heeee;
    LUT4 i21442_3_lut_4_lut (.A(\operand_1_x[2] ), .B(\operand_1_x[3] ), 
         .C(fill_value), .D(n93), .Z(n221)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i21442_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i21444_3_lut_4_lut (.A(\operand_1_x[2] ), .B(\operand_1_x[3] ), 
         .C(fill_value), .D(n94), .Z(n222)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i21444_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i21420_2_lut_rep_394 (.A(\operand_1_x[1] ), .B(\operand_1_x[2] ), 
         .Z(n41481)) /* synthesis lut_function=(A+(B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i21420_2_lut_rep_394.init = 16'heeee;
    LUT4 i21445_2_lut_rep_353_3_lut (.A(\operand_1_x[1] ), .B(\operand_1_x[2] ), 
         .C(\operand_1_x[3] ), .Z(n41440)) /* synthesis lut_function=(A+(B+(C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i21445_2_lut_rep_353_3_lut.init = 16'hfefe;
    LUT4 i21421_3_lut_4_lut (.A(\operand_1_x[1] ), .B(\operand_1_x[2] ), 
         .C(fill_value), .D(n31), .Z(n159)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i21421_3_lut_4_lut.init = 16'hf1e0;
    LUT4 i21415_2_lut_rep_395 (.A(\operand_1_x[0] ), .B(\operand_1_x[1] ), 
         .Z(n41482)) /* synthesis lut_function=(A+(B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i21415_2_lut_rep_395.init = 16'heeee;
    LUT4 i21422_2_lut_rep_354_3_lut (.A(\operand_1_x[0] ), .B(\operand_1_x[1] ), 
         .C(\operand_1_x[2] ), .Z(n41441)) /* synthesis lut_function=(A+(B+(C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i21422_2_lut_rep_354_3_lut.init = 16'hfefe;
    LUT4 i21447_2_lut_rep_327_3_lut_4_lut (.A(\operand_1_x[0] ), .B(\operand_1_x[1] ), 
         .C(\operand_1_x[3] ), .D(\operand_1_x[2] ), .Z(n41414)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i21447_2_lut_rep_327_3_lut_4_lut.init = 16'hfffe;
    LUT4 i21416_3_lut_4_lut (.A(\operand_1_x[0] ), .B(\operand_1_x[1] ), 
         .C(fill_value), .D(right_shift_operand[31]), .Z(n96)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(149[38:107])
    defparam i21416_3_lut_4_lut.init = 16'hf1e0;
    FD1P3AX right_shift_result_i0_i28 (.D(left_shift_result_31__N_2188[28]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i28.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i27 (.D(left_shift_result_31__N_2188[27]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i27.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i26 (.D(left_shift_result_31__N_2188[26]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[5])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i26.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i25 (.D(left_shift_result_31__N_2188[25]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[6])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i25.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i24 (.D(left_shift_result_31__N_2188[24]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[7])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i24.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i23 (.D(left_shift_result_31__N_2188[23]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[8])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i23.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i22 (.D(left_shift_result_31__N_2188[22]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[9])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i22.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i21 (.D(left_shift_result_31__N_2188[21]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[10])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i21.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i20 (.D(left_shift_result_31__N_2188[20]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[11])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i20.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i19 (.D(left_shift_result_31__N_2188[19]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[12])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i19.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i18 (.D(left_shift_result_31__N_2188[18]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[13])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i18.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i17 (.D(left_shift_result_31__N_2188[17]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[14])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i17.GSR = "ENABLED";
    PFUMX i37226 (.BLUT(n39778), .ALUT(n39779), .C0(\operand_1_x[4] ), 
          .Z(left_shift_result_31__N_2188[9]));
    FD1P3AX right_shift_result_i0_i16 (.D(left_shift_result_31__N_2188[16]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[15])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i16.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i15 (.D(left_shift_result_31__N_2188[15]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[16])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i15.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i14 (.D(left_shift_result_31__N_2188[14]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[17])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i14.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i13 (.D(left_shift_result_31__N_2188[13]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[18])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i13.GSR = "ENABLED";
    FD1P3AX right_shift_result_i0_i12 (.D(left_shift_result_31__N_2188[12]), 
            .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), .Q(left_shift_result[19])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=14, LSE_RCOL=6, LSE_LLINE=1071, LSE_RLINE=1082 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_shifter.v(146[5] 152[8])
    defparam right_shift_result_i0_i12.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module lm32_multiplier
//

module lm32_multiplier (GND_net, muliplicand, operand_1_x, multiplier_result_w, 
            w_clk_cpu, n41428, store_m, LM32D_CYC_O, n41512, w_clk_cpu_enable_623, 
            n46, reset_exception, n22524, \size_x[1] , \condition_x[0] , 
            n26122, n41513, data_bus_error_exception, memop_pc_w_31__N_1219, 
            w_clk_cpu_enable_972, w_clk_cpu_enable_984, n26142, \bypass_data_0[1] , 
            w_clk_cpu_enable_711, \bypass_data_0[0] , \d_result_0[31] , 
            \d_result_0[30] , \d_result_0[29] , \d_result_0[28] , \d_result_0[27] , 
            \d_result_0[26] , \d_result_0[25] , \d_result_0[24] , \d_result_0[23] , 
            \d_result_0[22] , \d_result_0[21] , \d_result_0[20] , \d_result_0[19] , 
            \d_result_0[18] , \d_result_0[17] , \d_result_0[16] , \d_result_0[15] , 
            \d_result_0[14] , \d_result_0[13] , \d_result_0[12] , \d_result_0[11] , 
            \d_result_0[10] , \d_result_0[9] , \d_result_0[8] , \d_result_0[7] , 
            \d_result_0[6] , \d_result_0[5] , \d_result_0[4] , \d_result_0[3] , 
            \d_result_0[2] ) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output [31:0]muliplicand;
    input [31:0]operand_1_x;
    output [31:0]multiplier_result_w;
    input w_clk_cpu;
    input n41428;
    input store_m;
    input LM32D_CYC_O;
    input n41512;
    output w_clk_cpu_enable_623;
    output n46;
    input reset_exception;
    output n22524;
    input \size_x[1] ;
    input \condition_x[0] ;
    output n26122;
    input n41513;
    input data_bus_error_exception;
    output memop_pc_w_31__N_1219;
    input w_clk_cpu_enable_972;
    input w_clk_cpu_enable_984;
    input n26142;
    input \bypass_data_0[1] ;
    input w_clk_cpu_enable_711;
    input \bypass_data_0[0] ;
    input \d_result_0[31] ;
    input \d_result_0[30] ;
    input \d_result_0[29] ;
    input \d_result_0[28] ;
    input \d_result_0[27] ;
    input \d_result_0[26] ;
    input \d_result_0[25] ;
    input \d_result_0[24] ;
    input \d_result_0[23] ;
    input \d_result_0[22] ;
    input \d_result_0[21] ;
    input \d_result_0[20] ;
    input \d_result_0[19] ;
    input \d_result_0[18] ;
    input \d_result_0[17] ;
    input \d_result_0[16] ;
    input \d_result_0[15] ;
    input \d_result_0[14] ;
    input \d_result_0[13] ;
    input \d_result_0[12] ;
    input \d_result_0[11] ;
    input \d_result_0[10] ;
    input \d_result_0[9] ;
    input \d_result_0[8] ;
    input \d_result_0[7] ;
    input \d_result_0[6] ;
    input \d_result_0[5] ;
    input \d_result_0[4] ;
    input \d_result_0[3] ;
    input \d_result_0[2] ;
    
    wire w_clk_cpu /* synthesis SET_AS_NETWORK=w_clk_cpu, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(22[6:15])
    
    wire mult_32u_32u_0_cin_lr_0, mult_32u_32u_0_pp_15_30, mult_32u_32u_0_pp_14_28, 
        mult_32u_32u_0_pp_13_26, mult_32u_32u_0_pp_12_24, mult_32u_32u_0_pp_11_22, 
        mult_32u_32u_0_pp_10_20, mult_32u_32u_0_pp_9_18, mult_32u_32u_0_pp_8_16, 
        mult_32u_32u_0_pp_7_14, mult_32u_32u_0_pp_6_12, mult_32u_32u_0_pp_5_10, 
        mult_32u_32u_0_pp_15_32, mult_32u_32u_0_pp_15_31, mult_32u_32u_0_cin_lr_30, 
        mult_32u_32u_0_pp_14_32, mult_32u_32u_0_pp_14_31, mco_210, mult_32u_32u_0_pp_14_30, 
        mult_32u_32u_0_pp_14_29, mult_32u_32u_0_cin_lr_28, co_mult_32u_32u_0_13_4, 
        s_mult_32u_32u_0_11_31, s_mult_32u_32u_0_11_32, s_mult_32u_32u_0_10_31, 
        s_mult_32u_32u_0_10_32, s_mult_32u_32u_0_13_31, s_mult_32u_32u_0_13_32, 
        co_mult_32u_32u_0_13_3, s_mult_32u_32u_0_11_29, s_mult_32u_32u_0_11_30, 
        s_mult_32u_32u_0_10_29, s_mult_32u_32u_0_10_30, s_mult_32u_32u_0_13_29, 
        s_mult_32u_32u_0_13_30, co_mult_32u_32u_0_13_2, s_mult_32u_32u_0_6_27, 
        s_mult_32u_32u_0_11_28, s_mult_32u_32u_0_10_27, s_mult_32u_32u_0_10_28, 
        s_mult_32u_32u_0_13_27, s_mult_32u_32u_0_13_28;
    wire [31:0]product;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(92[22:29])
    
    wire co_mult_32u_32u_0_13_1, s_mult_32u_32u_0_6_26, s_mult_32u_32u_0_10_25, 
        s_mult_32u_32u_0_10_26, s_mult_32u_32u_0_13_25, s_mult_32u_32u_0_13_26, 
        mult_32u_32u_0_pp_12_25, mult_32u_32u_0_pp_13_32, mult_32u_32u_0_pp_13_31, 
        mco_196, mult_32u_32u_0_pp_13_30, mult_32u_32u_0_pp_13_29, mco_195, 
        mult_32u_32u_0_pp_13_28, mult_32u_32u_0_pp_13_27, mult_32u_32u_0_cin_lr_26, 
        mult_32u_32u_0_pp_12_32, mult_32u_32u_0_pp_12_31, mco_182, mult_32u_32u_0_pp_12_30, 
        mult_32u_32u_0_pp_12_29, mco_181, mult_32u_32u_0_pp_12_28, mult_32u_32u_0_pp_12_27, 
        mco_180, mult_32u_32u_0_pp_12_26, mult_32u_32u_0_cin_lr_24, mult_32u_32u_0_pp_11_32, 
        mult_32u_32u_0_pp_11_31, mco_168, mult_32u_32u_0_pp_11_30, mult_32u_32u_0_pp_11_29, 
        mco_167, mult_32u_32u_0_pp_11_28, mult_32u_32u_0_pp_11_27, mco_166, 
        mult_32u_32u_0_pp_11_26, mult_32u_32u_0_pp_11_25, mco_165, mult_32u_32u_0_pp_11_24, 
        mult_32u_32u_0_pp_11_23, mult_32u_32u_0_cin_lr_22, mult_32u_32u_0_pp_10_32, 
        mult_32u_32u_0_pp_10_31, mco_154, mult_32u_32u_0_pp_10_30, mult_32u_32u_0_pp_10_29, 
        mco_153, mult_32u_32u_0_pp_10_28, mult_32u_32u_0_pp_10_27, mco_152, 
        mult_32u_32u_0_pp_10_26, mult_32u_32u_0_pp_10_25, mco_151, mult_32u_32u_0_pp_10_24, 
        mult_32u_32u_0_pp_10_23, mco_150, mult_32u_32u_0_pp_10_22, mult_32u_32u_0_pp_10_21, 
        mult_32u_32u_0_cin_lr_20, mult_32u_32u_0_pp_9_32, mult_32u_32u_0_pp_9_31, 
        mco_140, mult_32u_32u_0_pp_9_30, mult_32u_32u_0_pp_9_29, mco_139, 
        s_mult_32u_32u_0_10_24, s_mult_32u_32u_0_13_24, mult_32u_32u_0_pp_9_28, 
        mult_32u_32u_0_pp_9_27, mco_138, mult_32u_32u_0_pp_9_26, mult_32u_32u_0_pp_9_25, 
        mco_137, mult_32u_32u_0_pp_9_24, mult_32u_32u_0_pp_9_23, mco_136, 
        mult_32u_32u_0_pp_9_22, mult_32u_32u_0_pp_9_21, mco_135, mult_32u_32u_0_pp_9_20, 
        mult_32u_32u_0_pp_9_19, mult_32u_32u_0_cin_lr_18, mult_32u_32u_0_pp_8_32, 
        mult_32u_32u_0_pp_8_31, mco_126, mult_32u_32u_0_pp_8_30, mult_32u_32u_0_pp_8_29, 
        mco_125, mult_32u_32u_0_pp_8_28, mult_32u_32u_0_pp_8_27, mco_124, 
        mult_32u_32u_0_pp_8_26, mult_32u_32u_0_pp_8_25, mco_123, mult_32u_32u_0_pp_8_24, 
        mult_32u_32u_0_pp_8_23, mco_122, mult_32u_32u_0_pp_8_22, mult_32u_32u_0_pp_8_21, 
        mco_121, mult_32u_32u_0_pp_8_20, mult_32u_32u_0_pp_8_19, mco_120, 
        mult_32u_32u_0_pp_8_18, mult_32u_32u_0_pp_8_17, mult_32u_32u_0_cin_lr_16, 
        mult_32u_32u_0_pp_7_32, mult_32u_32u_0_pp_7_31, mco_112, mult_32u_32u_0_pp_7_30, 
        mult_32u_32u_0_pp_7_29, mco_111, mult_32u_32u_0_pp_7_28, mult_32u_32u_0_pp_7_27, 
        mco_110, mult_32u_32u_0_pp_7_26, mult_32u_32u_0_pp_7_25, mco_109, 
        mult_32u_32u_0_pp_7_24, mult_32u_32u_0_pp_7_23, mco_108, mult_32u_32u_0_pp_7_22, 
        mult_32u_32u_0_pp_7_21, mco_107, mult_32u_32u_0_pp_7_20, mult_32u_32u_0_pp_7_19, 
        mco_106, mult_32u_32u_0_pp_7_18, mult_32u_32u_0_pp_7_17, mco_105, 
        mult_32u_32u_0_pp_7_16, mult_32u_32u_0_pp_7_15, mult_32u_32u_0_cin_lr_14, 
        mult_32u_32u_0_pp_6_32, mult_32u_32u_0_pp_6_31, mco_98, mult_32u_32u_0_pp_6_30, 
        mult_32u_32u_0_pp_6_29, mco_97, mult_32u_32u_0_pp_6_28, mult_32u_32u_0_pp_6_27, 
        mco_96, mult_32u_32u_0_pp_6_26, mult_32u_32u_0_pp_6_25, mco_95, 
        mult_32u_32u_0_pp_6_24, mult_32u_32u_0_pp_6_23, mco_94, mult_32u_32u_0_pp_6_22, 
        mult_32u_32u_0_pp_6_21, mco_93, mult_32u_32u_0_pp_6_20, mult_32u_32u_0_pp_6_19, 
        mco_92, mult_32u_32u_0_pp_6_18, mult_32u_32u_0_pp_6_17, mco_91, 
        mult_32u_32u_0_pp_6_16, mult_32u_32u_0_pp_6_15, mco_90, mult_32u_32u_0_pp_6_14, 
        mult_32u_32u_0_pp_6_13, mult_32u_32u_0_cin_lr_12, mult_32u_32u_0_pp_5_32, 
        mult_32u_32u_0_pp_5_31, mco_84, mult_32u_32u_0_pp_5_30, mult_32u_32u_0_pp_5_29, 
        mco_83, mult_32u_32u_0_pp_5_28, mult_32u_32u_0_pp_5_27, mco_82, 
        mult_32u_32u_0_pp_5_26, mult_32u_32u_0_pp_5_25, mco_81, mult_32u_32u_0_pp_5_24, 
        mult_32u_32u_0_pp_5_23, mco_80, mult_32u_32u_0_pp_5_22, mult_32u_32u_0_pp_5_21, 
        mco_79, mult_32u_32u_0_pp_5_20, mult_32u_32u_0_pp_5_19, mco_78, 
        mult_32u_32u_0_pp_5_18, mult_32u_32u_0_pp_5_17, mco_77, mult_32u_32u_0_pp_5_16, 
        mult_32u_32u_0_pp_5_15, mco_76, mult_32u_32u_0_pp_5_14, mult_32u_32u_0_pp_5_13, 
        mco_75, mult_32u_32u_0_pp_5_12, mult_32u_32u_0_pp_5_11, mult_32u_32u_0_cin_lr_10, 
        co_mult_32u_32u_0_6_1, mult_32u_32u_0_pp_4_32, mult_32u_32u_0_pp_4_31, 
        mco_70, mult_32u_32u_0_pp_4_30, mult_32u_32u_0_pp_4_29, mco_69, 
        mult_32u_32u_0_pp_4_28, mult_32u_32u_0_pp_4_27, mco_68, mult_32u_32u_0_pp_4_26, 
        mult_32u_32u_0_pp_4_25, mco_67, mult_32u_32u_0_pp_4_24, mult_32u_32u_0_pp_4_23, 
        mco_66, mult_32u_32u_0_pp_4_22, mult_32u_32u_0_pp_4_21, mco_65, 
        mult_32u_32u_0_pp_4_20, mult_32u_32u_0_pp_4_19, mco_64, mult_32u_32u_0_pp_4_18, 
        mult_32u_32u_0_pp_4_17, mco_63, mult_32u_32u_0_pp_4_16, mult_32u_32u_0_pp_4_15, 
        mco_62, mult_32u_32u_0_pp_4_14, mult_32u_32u_0_pp_4_13, mco_61, 
        mult_32u_32u_0_pp_4_12, mult_32u_32u_0_pp_4_11, mco_60, mult_32u_32u_0_pp_4_10, 
        mult_32u_32u_0_pp_4_9, mult_32u_32u_0_cin_lr_8, mult_32u_32u_0_pp_3_32, 
        mult_32u_32u_0_pp_3_31, mco_56, mult_32u_32u_0_pp_3_30, mult_32u_32u_0_pp_3_29, 
        mco_55, mult_32u_32u_0_pp_3_28, mult_32u_32u_0_pp_3_27, mco_54, 
        mult_32u_32u_0_pp_3_26, mult_32u_32u_0_pp_3_25, mco_53, mult_32u_32u_0_pp_3_24, 
        mult_32u_32u_0_pp_3_23, mco_52, mult_32u_32u_0_pp_3_22, mult_32u_32u_0_pp_3_21, 
        mco_51, mult_32u_32u_0_pp_3_20, mult_32u_32u_0_pp_3_19, mco_50, 
        mult_32u_32u_0_pp_3_18, mult_32u_32u_0_pp_3_17, mco_49, mult_32u_32u_0_pp_3_16, 
        mult_32u_32u_0_pp_3_15, mco_48, mult_32u_32u_0_pp_3_14, mult_32u_32u_0_pp_3_13, 
        mco_47, mult_32u_32u_0_pp_3_12, mult_32u_32u_0_pp_3_11, mco_46, 
        mult_32u_32u_0_pp_3_10, mult_32u_32u_0_pp_3_9, mco_45, mult_32u_32u_0_pp_3_8, 
        mult_32u_32u_0_pp_3_7, mult_32u_32u_0_cin_lr_6, mult_32u_32u_0_pp_2_32, 
        mult_32u_32u_0_pp_2_31, mco_42, mult_32u_32u_0_pp_2_30, mult_32u_32u_0_pp_2_29, 
        mco_41, mult_32u_32u_0_pp_2_28, mult_32u_32u_0_pp_2_27, mco_40, 
        mult_32u_32u_0_pp_2_26, mult_32u_32u_0_pp_2_25, mco_39, mult_32u_32u_0_pp_2_24, 
        mult_32u_32u_0_pp_2_23, mco_38, mult_32u_32u_0_pp_2_22, mult_32u_32u_0_pp_2_21, 
        mco_37, mult_32u_32u_0_pp_2_20, mult_32u_32u_0_pp_2_19, mco_36, 
        mult_32u_32u_0_pp_2_18, mult_32u_32u_0_pp_2_17, mco_35, mult_32u_32u_0_pp_2_16, 
        mult_32u_32u_0_pp_2_15, mco_34, mult_32u_32u_0_pp_2_14, mult_32u_32u_0_pp_2_13, 
        mco_33, mult_32u_32u_0_pp_2_12, mult_32u_32u_0_pp_2_11, mco_32, 
        mult_32u_32u_0_pp_2_10, mult_32u_32u_0_pp_2_9, mco_31, mult_32u_32u_0_pp_2_8, 
        mult_32u_32u_0_pp_2_7, mco_30, mult_32u_32u_0_pp_2_6, mult_32u_32u_0_pp_2_5, 
        mult_32u_32u_0_cin_lr_4, mult_32u_32u_0_pp_1_32, mult_32u_32u_0_pp_1_31, 
        mco_28, mult_32u_32u_0_pp_1_30, mult_32u_32u_0_pp_1_29, mco_27, 
        mult_32u_32u_0_pp_1_28, mult_32u_32u_0_pp_1_27, mco_26, mult_32u_32u_0_pp_1_26, 
        mult_32u_32u_0_pp_1_25, mco_25, mult_32u_32u_0_pp_1_24, mult_32u_32u_0_pp_1_23, 
        mco_24, mult_32u_32u_0_pp_1_22, mult_32u_32u_0_pp_1_21, mco_23, 
        mult_32u_32u_0_pp_1_20, mult_32u_32u_0_pp_1_19, mco_22, mult_32u_32u_0_pp_1_18, 
        mult_32u_32u_0_pp_1_17, mco_21, mult_32u_32u_0_pp_1_16, mult_32u_32u_0_pp_1_15, 
        mco_20, mult_32u_32u_0_pp_1_14, mult_32u_32u_0_pp_1_13, mco_19, 
        mult_32u_32u_0_pp_1_12, mult_32u_32u_0_pp_1_11, mco_18, mult_32u_32u_0_pp_1_10, 
        mult_32u_32u_0_pp_1_9, mco_17, mult_32u_32u_0_pp_1_8, mult_32u_32u_0_pp_1_7, 
        mco_16, mult_32u_32u_0_pp_1_6, mult_32u_32u_0_pp_1_5, mco_15, 
        co_mult_32u_32u_0_4_7, s_mult_32u_32u_0_4_31, s_mult_32u_32u_0_4_32, 
        mult_32u_32u_0_pp_1_4, mult_32u_32u_0_pp_1_3, mult_32u_32u_0_cin_lr_2, 
        mult_32u_32u_0_pp_0_32, mult_32u_32u_0_pp_0_31, mco_14, co_mult_32u_32u_0_12_12, 
        s_mult_32u_32u_0_9_31, s_mult_32u_32u_0_9_32, s_mult_32u_32u_0_8_31, 
        s_mult_32u_32u_0_8_32, s_mult_32u_32u_0_12_31, s_mult_32u_32u_0_12_32, 
        mult_32u_32u_0_pp_0_30, mult_32u_32u_0_pp_0_29, mco_13, mult_32u_32u_0_pp_0_28, 
        mult_32u_32u_0_pp_0_27, mco_12, co_mult_32u_32u_0_12_11, s_mult_32u_32u_0_9_29, 
        s_mult_32u_32u_0_9_30, s_mult_32u_32u_0_8_29, s_mult_32u_32u_0_8_30, 
        s_mult_32u_32u_0_12_29, s_mult_32u_32u_0_12_30, co_mult_32u_32u_0_12_10, 
        s_mult_32u_32u_0_9_27, s_mult_32u_32u_0_9_28, s_mult_32u_32u_0_8_27, 
        s_mult_32u_32u_0_8_28, s_mult_32u_32u_0_12_27, s_mult_32u_32u_0_12_28, 
        co_mult_32u_32u_0_4_6, s_mult_32u_32u_0_4_29, s_mult_32u_32u_0_4_30, 
        co_mult_32u_32u_0_5_1, s_mult_32u_32u_0_5_22, mult_32u_32u_0_pp_0_26, 
        mult_32u_32u_0_pp_0_25, mco_11, co_mult_32u_32u_0_12_9, s_mult_32u_32u_0_9_25, 
        s_mult_32u_32u_0_9_26, s_mult_32u_32u_0_8_25, s_mult_32u_32u_0_8_26, 
        s_mult_32u_32u_0_12_25, s_mult_32u_32u_0_12_26, co_mult_32u_32u_0_12_8, 
        s_mult_32u_32u_0_9_23, s_mult_32u_32u_0_9_24, s_mult_32u_32u_0_8_23, 
        s_mult_32u_32u_0_8_24, s_mult_32u_32u_0_12_23, s_mult_32u_32u_0_12_24, 
        co_mult_32u_32u_0_4_5, s_mult_32u_32u_0_4_27, s_mult_32u_32u_0_4_28, 
        co_mult_32u_32u_0_4_4, s_mult_32u_32u_0_4_25, s_mult_32u_32u_0_4_26, 
        co_mult_32u_32u_0_12_7, s_mult_32u_32u_0_9_21, s_mult_32u_32u_0_9_22, 
        s_mult_32u_32u_0_8_21, s_mult_32u_32u_0_8_22, s_mult_32u_32u_0_12_21, 
        s_mult_32u_32u_0_12_22, co_mult_32u_32u_0_4_3, s_mult_32u_32u_0_4_23, 
        s_mult_32u_32u_0_4_24, co_mult_32u_32u_0_4_2, s_mult_32u_32u_0_4_21, 
        s_mult_32u_32u_0_4_22, co_mult_32u_32u_0_4_1, s_mult_32u_32u_0_4_20, 
        s_mult_32u_32u_0_4_19, co_mult_32u_32u_0_12_6, s_mult_32u_32u_0_9_19, 
        s_mult_32u_32u_0_9_20, s_mult_32u_32u_0_8_19, s_mult_32u_32u_0_8_20, 
        s_mult_32u_32u_0_12_19, s_mult_32u_32u_0_12_20, co_mult_32u_32u_0_12_5, 
        s_mult_32u_32u_0_9_17, s_mult_32u_32u_0_9_18, s_mult_32u_32u_0_8_17, 
        s_mult_32u_32u_0_8_18, s_mult_32u_32u_0_12_17, s_mult_32u_32u_0_12_18, 
        s_mult_32u_32u_0_4_18, mult_32u_32u_0_pp_0_24, mult_32u_32u_0_pp_0_23, 
        mco_10;
    wire [63:0]product_31__N_2324;
    
    wire co_mult_32u_32u_0_12_4, s_mult_32u_32u_0_9_15, s_mult_32u_32u_0_9_16, 
        s_mult_32u_32u_0_8_15, s_mult_32u_32u_0_8_16, s_mult_32u_32u_0_12_16, 
        mult_32u_32u_0_pp_0_22, mult_32u_32u_0_pp_0_21, mco_9, mult_32u_32u_0_pp_0_20, 
        mult_32u_32u_0_pp_0_19, mco_8, mult_32u_32u_0_pp_0_18, mult_32u_32u_0_pp_0_17, 
        mco_7, mult_32u_32u_0_pp_0_16, mult_32u_32u_0_pp_0_15, mco_6, 
        mult_32u_32u_0_pp_0_14, mult_32u_32u_0_pp_0_13, mco_5, co_mult_32u_32u_0_12_3, 
        s_mult_32u_32u_0_9_13, s_mult_32u_32u_0_9_14, s_mult_32u_32u_0_8_13, 
        s_mult_32u_32u_0_8_14, mult_32u_32u_0_pp_0_12, mult_32u_32u_0_pp_0_11, 
        mco_4, co_mult_32u_32u_0_12_2, s_mult_32u_32u_0_2_11, s_mult_32u_32u_0_9_12, 
        s_mult_32u_32u_0_8_11, s_mult_32u_32u_0_8_12, mult_32u_32u_0_pp_0_10, 
        mult_32u_32u_0_pp_0_9, mco_3, co_mult_32u_32u_0_12_1, s_mult_32u_32u_0_2_10, 
        s_mult_32u_32u_0_8_9, s_mult_32u_32u_0_8_10, mult_32u_32u_0_pp_0_8, 
        mult_32u_32u_0_pp_0_7, mco_2, mult_32u_32u_0_pp_4_8, s_mult_32u_32u_0_8_8, 
        mult_32u_32u_0_pp_0_6, mult_32u_32u_0_pp_0_5, mco_1, mult_32u_32u_0_pp_0_4, 
        mult_32u_32u_0_pp_0_3, mco, mult_32u_32u_0_pp_0_2, co_t_mult_32u_32u_0_14_8, 
        co_t_mult_32u_32u_0_14_7, co_t_mult_32u_32u_0_14_6, co_t_mult_32u_32u_0_14_5, 
        co_t_mult_32u_32u_0_14_4, s_mult_32u_32u_0_10_23, co_t_mult_32u_32u_0_14_3, 
        s_mult_32u_32u_0_10_21, s_mult_32u_32u_0_10_22, co_t_mult_32u_32u_0_14_2, 
        s_mult_32u_32u_0_10_20, co_t_mult_32u_32u_0_14_1, co_mult_32u_32u_0_3_9, 
        s_mult_32u_32u_0_3_31, s_mult_32u_32u_0_3_32, co_mult_32u_32u_0_3_8, 
        s_mult_32u_32u_0_3_29, s_mult_32u_32u_0_3_30, co_mult_32u_32u_0_3_7, 
        s_mult_32u_32u_0_3_27, s_mult_32u_32u_0_3_28, co_mult_32u_32u_0_3_6, 
        s_mult_32u_32u_0_3_25, s_mult_32u_32u_0_3_26, co_mult_32u_32u_0_3_5, 
        s_mult_32u_32u_0_3_23, s_mult_32u_32u_0_3_24, co_mult_32u_32u_0_3_4, 
        s_mult_32u_32u_0_3_21, s_mult_32u_32u_0_3_22, co_mult_32u_32u_0_3_3, 
        s_mult_32u_32u_0_3_19, s_mult_32u_32u_0_3_20, co_mult_32u_32u_0_3_2, 
        s_mult_32u_32u_0_3_17, s_mult_32u_32u_0_3_18, co_mult_32u_32u_0_3_1, 
        s_mult_32u_32u_0_3_15, s_mult_32u_32u_0_3_16, s_mult_32u_32u_0_3_14, 
        co_mult_32u_32u_0_11_2, s_mult_32u_32u_0_7_31, s_mult_32u_32u_0_7_32, 
        s_mult_32u_32u_0_6_31, s_mult_32u_32u_0_6_32, co_mult_32u_32u_0_11_1, 
        s_mult_32u_32u_0_7_30, s_mult_32u_32u_0_6_29, s_mult_32u_32u_0_6_30, 
        co_mult_32u_32u_0_2_11, s_mult_32u_32u_0_2_31, s_mult_32u_32u_0_2_32, 
        s_mult_32u_32u_0_6_28, co_mult_32u_32u_0_2_10, s_mult_32u_32u_0_2_29, 
        s_mult_32u_32u_0_2_30, co_mult_32u_32u_0_2_9, s_mult_32u_32u_0_2_27, 
        s_mult_32u_32u_0_2_28, co_mult_32u_32u_0_2_8, s_mult_32u_32u_0_2_25, 
        s_mult_32u_32u_0_2_26, co_mult_32u_32u_0_2_7, s_mult_32u_32u_0_2_23, 
        s_mult_32u_32u_0_2_24, co_mult_32u_32u_0_2_6, s_mult_32u_32u_0_2_21, 
        s_mult_32u_32u_0_2_22, co_mult_32u_32u_0_2_5, s_mult_32u_32u_0_2_19, 
        s_mult_32u_32u_0_2_20, co_mult_32u_32u_0_2_4, s_mult_32u_32u_0_2_17, 
        s_mult_32u_32u_0_2_18, co_mult_32u_32u_0_2_3, s_mult_32u_32u_0_2_15, 
        s_mult_32u_32u_0_2_16, co_mult_32u_32u_0_2_2, s_mult_32u_32u_0_2_13, 
        s_mult_32u_32u_0_2_14, co_mult_32u_32u_0_10_6, s_mult_32u_32u_0_5_31, 
        s_mult_32u_32u_0_5_32, co_mult_32u_32u_0_10_5, s_mult_32u_32u_0_5_29, 
        s_mult_32u_32u_0_5_30, co_mult_32u_32u_0_10_4, s_mult_32u_32u_0_5_27, 
        s_mult_32u_32u_0_5_28, co_mult_32u_32u_0_2_1, s_mult_32u_32u_0_2_12, 
        co_mult_32u_32u_0_10_3, s_mult_32u_32u_0_5_25, s_mult_32u_32u_0_5_26, 
        co_mult_32u_32u_0_10_2, s_mult_32u_32u_0_5_23, s_mult_32u_32u_0_5_24, 
        co_mult_32u_32u_0_10_1, co_mult_32u_32u_0_1_13, s_mult_32u_32u_0_1_31, 
        s_mult_32u_32u_0_1_32, co_mult_32u_32u_0_1_12, s_mult_32u_32u_0_1_29, 
        s_mult_32u_32u_0_1_30, co_mult_32u_32u_0_1_11, s_mult_32u_32u_0_1_27, 
        s_mult_32u_32u_0_1_28, co_mult_32u_32u_0_1_10, s_mult_32u_32u_0_1_25, 
        s_mult_32u_32u_0_1_26, co_mult_32u_32u_0_1_9, s_mult_32u_32u_0_1_23, 
        s_mult_32u_32u_0_1_24, co_mult_32u_32u_0_1_8, s_mult_32u_32u_0_1_21, 
        s_mult_32u_32u_0_1_22, co_mult_32u_32u_0_1_7, s_mult_32u_32u_0_1_19, 
        s_mult_32u_32u_0_1_20, co_mult_32u_32u_0_9_10, co_mult_32u_32u_0_9_9, 
        co_mult_32u_32u_0_1_6, s_mult_32u_32u_0_1_17, s_mult_32u_32u_0_1_18, 
        co_mult_32u_32u_0_1_5, s_mult_32u_32u_0_1_15, s_mult_32u_32u_0_1_16, 
        co_mult_32u_32u_0_1_4, s_mult_32u_32u_0_1_13, s_mult_32u_32u_0_1_14, 
        co_mult_32u_32u_0_1_3, s_mult_32u_32u_0_1_11, s_mult_32u_32u_0_1_12, 
        co_mult_32u_32u_0_1_2, s_mult_32u_32u_0_1_9, s_mult_32u_32u_0_1_10, 
        co_mult_32u_32u_0_1_1, s_mult_32u_32u_0_1_7, s_mult_32u_32u_0_1_8, 
        mult_32u_32u_0_pp_3_6, s_mult_32u_32u_0_1_6, co_mult_32u_32u_0_9_8, 
        co_mult_32u_32u_0_9_7, co_mult_32u_32u_0_0_15, s_mult_32u_32u_0_0_31, 
        s_mult_32u_32u_0_0_32, co_mult_32u_32u_0_0_14, s_mult_32u_32u_0_0_29, 
        s_mult_32u_32u_0_0_30, co_mult_32u_32u_0_0_13, s_mult_32u_32u_0_0_27, 
        s_mult_32u_32u_0_0_28, co_mult_32u_32u_0_0_12, s_mult_32u_32u_0_0_25, 
        s_mult_32u_32u_0_0_26, co_mult_32u_32u_0_0_11, s_mult_32u_32u_0_0_23, 
        s_mult_32u_32u_0_0_24, co_mult_32u_32u_0_0_10, s_mult_32u_32u_0_0_21, 
        s_mult_32u_32u_0_0_22, co_mult_32u_32u_0_9_6, co_mult_32u_32u_0_0_9, 
        s_mult_32u_32u_0_0_19, s_mult_32u_32u_0_0_20, co_mult_32u_32u_0_0_8, 
        s_mult_32u_32u_0_0_17, s_mult_32u_32u_0_0_18, co_mult_32u_32u_0_9_5, 
        co_mult_32u_32u_0_0_7, s_mult_32u_32u_0_0_15, s_mult_32u_32u_0_0_16, 
        co_mult_32u_32u_0_9_4, co_mult_32u_32u_0_0_6, s_mult_32u_32u_0_0_13, 
        s_mult_32u_32u_0_0_14, co_mult_32u_32u_0_0_5, s_mult_32u_32u_0_0_11, 
        s_mult_32u_32u_0_0_12, co_mult_32u_32u_0_0_4, s_mult_32u_32u_0_0_9, 
        s_mult_32u_32u_0_0_10, co_mult_32u_32u_0_0_3, s_mult_32u_32u_0_0_7, 
        s_mult_32u_32u_0_0_8, co_mult_32u_32u_0_0_2, s_mult_32u_32u_0_0_5, 
        s_mult_32u_32u_0_0_6, co_mult_32u_32u_0_0_1, s_mult_32u_32u_0_0_4, 
        mult_32u_32u_0_pp_1_2, co_mult_32u_32u_0_9_3, co_mult_32u_32u_0_9_2, 
        co_mult_32u_32u_0_9_1, mult_32u_32u_0_pp_2_4, co_mult_32u_32u_0_8_14, 
        co_mult_32u_32u_0_8_13, co_mult_32u_32u_0_8_12, co_mult_32u_32u_0_8_11, 
        co_mult_32u_32u_0_8_10, co_mult_32u_32u_0_8_9, co_mult_32u_32u_0_8_8, 
        co_mult_32u_32u_0_8_7, co_mult_32u_32u_0_8_6, co_mult_32u_32u_0_8_5, 
        co_mult_32u_32u_0_8_4, co_mult_32u_32u_0_8_3, co_mult_32u_32u_0_8_2, 
        co_mult_32u_32u_0_8_1, co_mult_32u_32u_0_7_1, co_mult_32u_32u_0_5_5, 
        co_mult_32u_32u_0_5_4, co_mult_32u_32u_0_5_3, co_mult_32u_32u_0_5_2, 
        co_mult_32u_32u_0_6_3, co_mult_32u_32u_0_6_2;
    
    FADD2B mult_32u_32u_0_cin_lr_add_0 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_32u_32u_0_cin_lr_0)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    AND2 AND2_t0 (.A(muliplicand[0]), .B(operand_1_x[30]), .Z(mult_32u_32u_0_pp_15_30)) /* synthesis syn_instantiated=1 */ ;   // mult_32u_32u.v(1684[10:68])
    AND2 AND2_t1 (.A(muliplicand[0]), .B(operand_1_x[28]), .Z(mult_32u_32u_0_pp_14_28)) /* synthesis syn_instantiated=1 */ ;   // mult_32u_32u.v(1682[10:68])
    AND2 AND2_t2 (.A(muliplicand[0]), .B(operand_1_x[26]), .Z(mult_32u_32u_0_pp_13_26)) /* synthesis syn_instantiated=1 */ ;   // mult_32u_32u.v(1680[10:68])
    AND2 AND2_t3 (.A(muliplicand[0]), .B(operand_1_x[24]), .Z(mult_32u_32u_0_pp_12_24)) /* synthesis syn_instantiated=1 */ ;   // mult_32u_32u.v(1678[10:68])
    AND2 AND2_t4 (.A(muliplicand[0]), .B(operand_1_x[22]), .Z(mult_32u_32u_0_pp_11_22)) /* synthesis syn_instantiated=1 */ ;   // mult_32u_32u.v(1676[10:68])
    AND2 AND2_t5 (.A(muliplicand[0]), .B(operand_1_x[20]), .Z(mult_32u_32u_0_pp_10_20)) /* synthesis syn_instantiated=1 */ ;   // mult_32u_32u.v(1674[10:68])
    AND2 AND2_t6 (.A(muliplicand[0]), .B(operand_1_x[18]), .Z(mult_32u_32u_0_pp_9_18)) /* synthesis syn_instantiated=1 */ ;   // mult_32u_32u.v(1672[10:67])
    AND2 AND2_t7 (.A(muliplicand[0]), .B(operand_1_x[16]), .Z(mult_32u_32u_0_pp_8_16)) /* synthesis syn_instantiated=1 */ ;   // mult_32u_32u.v(1670[10:67])
    AND2 AND2_t8 (.A(muliplicand[0]), .B(operand_1_x[14]), .Z(mult_32u_32u_0_pp_7_14)) /* synthesis syn_instantiated=1 */ ;   // mult_32u_32u.v(1668[10:67])
    AND2 AND2_t9 (.A(muliplicand[0]), .B(operand_1_x[12]), .Z(mult_32u_32u_0_pp_6_12)) /* synthesis syn_instantiated=1 */ ;   // mult_32u_32u.v(1666[10:67])
    AND2 AND2_t10 (.A(muliplicand[0]), .B(operand_1_x[10]), .Z(mult_32u_32u_0_pp_5_10)) /* synthesis syn_instantiated=1 */ ;   // mult_32u_32u.v(1664[10:68])
    MULT2 mult_32u_32u_0_mult_30_0 (.A0(muliplicand[0]), .A1(muliplicand[1]), 
          .A2(muliplicand[1]), .A3(muliplicand[2]), .B0(operand_1_x[31]), 
          .B1(operand_1_x[30]), .B2(operand_1_x[31]), .B3(operand_1_x[30]), 
          .CI(mult_32u_32u_0_cin_lr_30), .P0(mult_32u_32u_0_pp_15_31), .P1(mult_32u_32u_0_pp_15_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_28_1 (.A0(muliplicand[2]), .A1(muliplicand[3]), 
          .A2(muliplicand[3]), .A3(muliplicand[4]), .B0(operand_1_x[29]), 
          .B1(operand_1_x[28]), .B2(operand_1_x[29]), .B3(operand_1_x[28]), 
          .CI(mco_210), .P0(mult_32u_32u_0_pp_14_31), .P1(mult_32u_32u_0_pp_14_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_28_0 (.A0(muliplicand[0]), .A1(muliplicand[1]), 
          .A2(muliplicand[1]), .A3(muliplicand[2]), .B0(operand_1_x[29]), 
          .B1(operand_1_x[28]), .B2(operand_1_x[29]), .B3(operand_1_x[28]), 
          .CI(mult_32u_32u_0_cin_lr_28), .CO(mco_210), .P0(mult_32u_32u_0_pp_14_29), 
          .P1(mult_32u_32u_0_pp_14_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_13_5 (.A0(s_mult_32u_32u_0_10_31), .A1(s_mult_32u_32u_0_10_32), 
           .B0(s_mult_32u_32u_0_11_31), .B1(s_mult_32u_32u_0_11_32), .CI(co_mult_32u_32u_0_13_4), 
           .S0(s_mult_32u_32u_0_13_31), .S1(s_mult_32u_32u_0_13_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_13_4 (.A0(s_mult_32u_32u_0_10_29), .A1(s_mult_32u_32u_0_10_30), 
           .B0(s_mult_32u_32u_0_11_29), .B1(s_mult_32u_32u_0_11_30), .CI(co_mult_32u_32u_0_13_3), 
           .COUT(co_mult_32u_32u_0_13_4), .S0(s_mult_32u_32u_0_13_29), .S1(s_mult_32u_32u_0_13_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_13_3 (.A0(s_mult_32u_32u_0_10_27), .A1(s_mult_32u_32u_0_10_28), 
           .B0(s_mult_32u_32u_0_6_27), .B1(s_mult_32u_32u_0_11_28), .CI(co_mult_32u_32u_0_13_2), 
           .COUT(co_mult_32u_32u_0_13_3), .S0(s_mult_32u_32u_0_13_27), .S1(s_mult_32u_32u_0_13_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1S3AX result_i26 (.D(product[26]), .CK(w_clk_cpu), .Q(multiplier_result_w[26])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i26.GSR = "ENABLED";
    FADD2B mult_32u_32u_0_add_13_2 (.A0(s_mult_32u_32u_0_10_25), .A1(s_mult_32u_32u_0_10_26), 
           .B0(mult_32u_32u_0_pp_12_25), .B1(s_mult_32u_32u_0_6_26), .CI(co_mult_32u_32u_0_13_1), 
           .COUT(co_mult_32u_32u_0_13_2), .S0(s_mult_32u_32u_0_13_25), .S1(s_mult_32u_32u_0_13_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_26_2 (.A0(muliplicand[4]), .A1(muliplicand[5]), 
          .A2(muliplicand[5]), .A3(muliplicand[6]), .B0(operand_1_x[27]), 
          .B1(operand_1_x[26]), .B2(operand_1_x[27]), .B3(operand_1_x[26]), 
          .CI(mco_196), .P0(mult_32u_32u_0_pp_13_31), .P1(mult_32u_32u_0_pp_13_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_26_1 (.A0(muliplicand[2]), .A1(muliplicand[3]), 
          .A2(muliplicand[3]), .A3(muliplicand[4]), .B0(operand_1_x[27]), 
          .B1(operand_1_x[26]), .B2(operand_1_x[27]), .B3(operand_1_x[26]), 
          .CI(mco_195), .CO(mco_196), .P0(mult_32u_32u_0_pp_13_29), .P1(mult_32u_32u_0_pp_13_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_26_0 (.A0(muliplicand[0]), .A1(muliplicand[1]), 
          .A2(muliplicand[1]), .A3(muliplicand[2]), .B0(operand_1_x[27]), 
          .B1(operand_1_x[26]), .B2(operand_1_x[27]), .B3(operand_1_x[26]), 
          .CI(mult_32u_32u_0_cin_lr_26), .CO(mco_195), .P0(mult_32u_32u_0_pp_13_27), 
          .P1(mult_32u_32u_0_pp_13_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_24_3 (.A0(muliplicand[6]), .A1(muliplicand[7]), 
          .A2(muliplicand[7]), .A3(muliplicand[8]), .B0(operand_1_x[25]), 
          .B1(operand_1_x[24]), .B2(operand_1_x[25]), .B3(operand_1_x[24]), 
          .CI(mco_182), .P0(mult_32u_32u_0_pp_12_31), .P1(mult_32u_32u_0_pp_12_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_24_2 (.A0(muliplicand[4]), .A1(muliplicand[5]), 
          .A2(muliplicand[5]), .A3(muliplicand[6]), .B0(operand_1_x[25]), 
          .B1(operand_1_x[24]), .B2(operand_1_x[25]), .B3(operand_1_x[24]), 
          .CI(mco_181), .CO(mco_182), .P0(mult_32u_32u_0_pp_12_29), .P1(mult_32u_32u_0_pp_12_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_24_1 (.A0(muliplicand[2]), .A1(muliplicand[3]), 
          .A2(muliplicand[3]), .A3(muliplicand[4]), .B0(operand_1_x[25]), 
          .B1(operand_1_x[24]), .B2(operand_1_x[25]), .B3(operand_1_x[24]), 
          .CI(mco_180), .CO(mco_181), .P0(mult_32u_32u_0_pp_12_27), .P1(mult_32u_32u_0_pp_12_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_24_0 (.A0(muliplicand[0]), .A1(muliplicand[1]), 
          .A2(muliplicand[1]), .A3(muliplicand[2]), .B0(operand_1_x[25]), 
          .B1(operand_1_x[24]), .B2(operand_1_x[25]), .B3(operand_1_x[24]), 
          .CI(mult_32u_32u_0_cin_lr_24), .CO(mco_180), .P0(mult_32u_32u_0_pp_12_25), 
          .P1(mult_32u_32u_0_pp_12_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_22_4 (.A0(muliplicand[8]), .A1(muliplicand[9]), 
          .A2(muliplicand[9]), .A3(muliplicand[10]), .B0(operand_1_x[23]), 
          .B1(operand_1_x[22]), .B2(operand_1_x[23]), .B3(operand_1_x[22]), 
          .CI(mco_168), .P0(mult_32u_32u_0_pp_11_31), .P1(mult_32u_32u_0_pp_11_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_22_3 (.A0(muliplicand[6]), .A1(muliplicand[7]), 
          .A2(muliplicand[7]), .A3(muliplicand[8]), .B0(operand_1_x[23]), 
          .B1(operand_1_x[22]), .B2(operand_1_x[23]), .B3(operand_1_x[22]), 
          .CI(mco_167), .CO(mco_168), .P0(mult_32u_32u_0_pp_11_29), .P1(mult_32u_32u_0_pp_11_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_22_2 (.A0(muliplicand[4]), .A1(muliplicand[5]), 
          .A2(muliplicand[5]), .A3(muliplicand[6]), .B0(operand_1_x[23]), 
          .B1(operand_1_x[22]), .B2(operand_1_x[23]), .B3(operand_1_x[22]), 
          .CI(mco_166), .CO(mco_167), .P0(mult_32u_32u_0_pp_11_27), .P1(mult_32u_32u_0_pp_11_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_22_1 (.A0(muliplicand[2]), .A1(muliplicand[3]), 
          .A2(muliplicand[3]), .A3(muliplicand[4]), .B0(operand_1_x[23]), 
          .B1(operand_1_x[22]), .B2(operand_1_x[23]), .B3(operand_1_x[22]), 
          .CI(mco_165), .CO(mco_166), .P0(mult_32u_32u_0_pp_11_25), .P1(mult_32u_32u_0_pp_11_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_22_0 (.A0(muliplicand[0]), .A1(muliplicand[1]), 
          .A2(muliplicand[1]), .A3(muliplicand[2]), .B0(operand_1_x[23]), 
          .B1(operand_1_x[22]), .B2(operand_1_x[23]), .B3(operand_1_x[22]), 
          .CI(mult_32u_32u_0_cin_lr_22), .CO(mco_165), .P0(mult_32u_32u_0_pp_11_23), 
          .P1(mult_32u_32u_0_pp_11_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_20_5 (.A0(muliplicand[10]), .A1(muliplicand[11]), 
          .A2(muliplicand[11]), .A3(muliplicand[12]), .B0(operand_1_x[21]), 
          .B1(operand_1_x[20]), .B2(operand_1_x[21]), .B3(operand_1_x[20]), 
          .CI(mco_154), .P0(mult_32u_32u_0_pp_10_31), .P1(mult_32u_32u_0_pp_10_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_20_4 (.A0(muliplicand[8]), .A1(muliplicand[9]), 
          .A2(muliplicand[9]), .A3(muliplicand[10]), .B0(operand_1_x[21]), 
          .B1(operand_1_x[20]), .B2(operand_1_x[21]), .B3(operand_1_x[20]), 
          .CI(mco_153), .CO(mco_154), .P0(mult_32u_32u_0_pp_10_29), .P1(mult_32u_32u_0_pp_10_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_20_3 (.A0(muliplicand[6]), .A1(muliplicand[7]), 
          .A2(muliplicand[7]), .A3(muliplicand[8]), .B0(operand_1_x[21]), 
          .B1(operand_1_x[20]), .B2(operand_1_x[21]), .B3(operand_1_x[20]), 
          .CI(mco_152), .CO(mco_153), .P0(mult_32u_32u_0_pp_10_27), .P1(mult_32u_32u_0_pp_10_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_20_2 (.A0(muliplicand[4]), .A1(muliplicand[5]), 
          .A2(muliplicand[5]), .A3(muliplicand[6]), .B0(operand_1_x[21]), 
          .B1(operand_1_x[20]), .B2(operand_1_x[21]), .B3(operand_1_x[20]), 
          .CI(mco_151), .CO(mco_152), .P0(mult_32u_32u_0_pp_10_25), .P1(mult_32u_32u_0_pp_10_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_20_1 (.A0(muliplicand[2]), .A1(muliplicand[3]), 
          .A2(muliplicand[3]), .A3(muliplicand[4]), .B0(operand_1_x[21]), 
          .B1(operand_1_x[20]), .B2(operand_1_x[21]), .B3(operand_1_x[20]), 
          .CI(mco_150), .CO(mco_151), .P0(mult_32u_32u_0_pp_10_23), .P1(mult_32u_32u_0_pp_10_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_20_0 (.A0(muliplicand[0]), .A1(muliplicand[1]), 
          .A2(muliplicand[1]), .A3(muliplicand[2]), .B0(operand_1_x[21]), 
          .B1(operand_1_x[20]), .B2(operand_1_x[21]), .B3(operand_1_x[20]), 
          .CI(mult_32u_32u_0_cin_lr_20), .CO(mco_150), .P0(mult_32u_32u_0_pp_10_21), 
          .P1(mult_32u_32u_0_pp_10_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1S3AX result_i25 (.D(product[25]), .CK(w_clk_cpu), .Q(multiplier_result_w[25])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i25.GSR = "ENABLED";
    FD1S3AX result_i24 (.D(product[24]), .CK(w_clk_cpu), .Q(multiplier_result_w[24])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i24.GSR = "ENABLED";
    FD1S3AX result_i23 (.D(product[23]), .CK(w_clk_cpu), .Q(multiplier_result_w[23])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i23.GSR = "ENABLED";
    MULT2 mult_32u_32u_0_mult_18_6 (.A0(muliplicand[12]), .A1(muliplicand[13]), 
          .A2(muliplicand[13]), .A3(muliplicand[14]), .B0(operand_1_x[19]), 
          .B1(operand_1_x[18]), .B2(operand_1_x[19]), .B3(operand_1_x[18]), 
          .CI(mco_140), .P0(mult_32u_32u_0_pp_9_31), .P1(mult_32u_32u_0_pp_9_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_18_5 (.A0(muliplicand[10]), .A1(muliplicand[11]), 
          .A2(muliplicand[11]), .A3(muliplicand[12]), .B0(operand_1_x[19]), 
          .B1(operand_1_x[18]), .B2(operand_1_x[19]), .B3(operand_1_x[18]), 
          .CI(mco_139), .CO(mco_140), .P0(mult_32u_32u_0_pp_9_29), .P1(mult_32u_32u_0_pp_9_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B Cadd_mult_32u_32u_0_13_1 (.A0(GND_net), .A1(s_mult_32u_32u_0_10_24), 
           .B0(GND_net), .B1(mult_32u_32u_0_pp_12_24), .CI(GND_net), .COUT(co_mult_32u_32u_0_13_1), 
           .S1(s_mult_32u_32u_0_13_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_18_4 (.A0(muliplicand[8]), .A1(muliplicand[9]), 
          .A2(muliplicand[9]), .A3(muliplicand[10]), .B0(operand_1_x[19]), 
          .B1(operand_1_x[18]), .B2(operand_1_x[19]), .B3(operand_1_x[18]), 
          .CI(mco_138), .CO(mco_139), .P0(mult_32u_32u_0_pp_9_27), .P1(mult_32u_32u_0_pp_9_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_18_3 (.A0(muliplicand[6]), .A1(muliplicand[7]), 
          .A2(muliplicand[7]), .A3(muliplicand[8]), .B0(operand_1_x[19]), 
          .B1(operand_1_x[18]), .B2(operand_1_x[19]), .B3(operand_1_x[18]), 
          .CI(mco_137), .CO(mco_138), .P0(mult_32u_32u_0_pp_9_25), .P1(mult_32u_32u_0_pp_9_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_18_2 (.A0(muliplicand[4]), .A1(muliplicand[5]), 
          .A2(muliplicand[5]), .A3(muliplicand[6]), .B0(operand_1_x[19]), 
          .B1(operand_1_x[18]), .B2(operand_1_x[19]), .B3(operand_1_x[18]), 
          .CI(mco_136), .CO(mco_137), .P0(mult_32u_32u_0_pp_9_23), .P1(mult_32u_32u_0_pp_9_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_18_1 (.A0(muliplicand[2]), .A1(muliplicand[3]), 
          .A2(muliplicand[3]), .A3(muliplicand[4]), .B0(operand_1_x[19]), 
          .B1(operand_1_x[18]), .B2(operand_1_x[19]), .B3(operand_1_x[18]), 
          .CI(mco_135), .CO(mco_136), .P0(mult_32u_32u_0_pp_9_21), .P1(mult_32u_32u_0_pp_9_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_18_0 (.A0(muliplicand[0]), .A1(muliplicand[1]), 
          .A2(muliplicand[1]), .A3(muliplicand[2]), .B0(operand_1_x[19]), 
          .B1(operand_1_x[18]), .B2(operand_1_x[19]), .B3(operand_1_x[18]), 
          .CI(mult_32u_32u_0_cin_lr_18), .CO(mco_135), .P0(mult_32u_32u_0_pp_9_19), 
          .P1(mult_32u_32u_0_pp_9_20)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_16_7 (.A0(muliplicand[14]), .A1(muliplicand[15]), 
          .A2(muliplicand[15]), .A3(muliplicand[16]), .B0(operand_1_x[17]), 
          .B1(operand_1_x[16]), .B2(operand_1_x[17]), .B3(operand_1_x[16]), 
          .CI(mco_126), .P0(mult_32u_32u_0_pp_8_31), .P1(mult_32u_32u_0_pp_8_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_16_6 (.A0(muliplicand[12]), .A1(muliplicand[13]), 
          .A2(muliplicand[13]), .A3(muliplicand[14]), .B0(operand_1_x[17]), 
          .B1(operand_1_x[16]), .B2(operand_1_x[17]), .B3(operand_1_x[16]), 
          .CI(mco_125), .CO(mco_126), .P0(mult_32u_32u_0_pp_8_29), .P1(mult_32u_32u_0_pp_8_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_16_5 (.A0(muliplicand[10]), .A1(muliplicand[11]), 
          .A2(muliplicand[11]), .A3(muliplicand[12]), .B0(operand_1_x[17]), 
          .B1(operand_1_x[16]), .B2(operand_1_x[17]), .B3(operand_1_x[16]), 
          .CI(mco_124), .CO(mco_125), .P0(mult_32u_32u_0_pp_8_27), .P1(mult_32u_32u_0_pp_8_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_16_4 (.A0(muliplicand[8]), .A1(muliplicand[9]), 
          .A2(muliplicand[9]), .A3(muliplicand[10]), .B0(operand_1_x[17]), 
          .B1(operand_1_x[16]), .B2(operand_1_x[17]), .B3(operand_1_x[16]), 
          .CI(mco_123), .CO(mco_124), .P0(mult_32u_32u_0_pp_8_25), .P1(mult_32u_32u_0_pp_8_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_16_3 (.A0(muliplicand[6]), .A1(muliplicand[7]), 
          .A2(muliplicand[7]), .A3(muliplicand[8]), .B0(operand_1_x[17]), 
          .B1(operand_1_x[16]), .B2(operand_1_x[17]), .B3(operand_1_x[16]), 
          .CI(mco_122), .CO(mco_123), .P0(mult_32u_32u_0_pp_8_23), .P1(mult_32u_32u_0_pp_8_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_16_2 (.A0(muliplicand[4]), .A1(muliplicand[5]), 
          .A2(muliplicand[5]), .A3(muliplicand[6]), .B0(operand_1_x[17]), 
          .B1(operand_1_x[16]), .B2(operand_1_x[17]), .B3(operand_1_x[16]), 
          .CI(mco_121), .CO(mco_122), .P0(mult_32u_32u_0_pp_8_21), .P1(mult_32u_32u_0_pp_8_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1S3AX result_i22 (.D(product[22]), .CK(w_clk_cpu), .Q(multiplier_result_w[22])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i22.GSR = "ENABLED";
    MULT2 mult_32u_32u_0_mult_16_1 (.A0(muliplicand[2]), .A1(muliplicand[3]), 
          .A2(muliplicand[3]), .A3(muliplicand[4]), .B0(operand_1_x[17]), 
          .B1(operand_1_x[16]), .B2(operand_1_x[17]), .B3(operand_1_x[16]), 
          .CI(mco_120), .CO(mco_121), .P0(mult_32u_32u_0_pp_8_19), .P1(mult_32u_32u_0_pp_8_20)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_16_0 (.A0(muliplicand[0]), .A1(muliplicand[1]), 
          .A2(muliplicand[1]), .A3(muliplicand[2]), .B0(operand_1_x[17]), 
          .B1(operand_1_x[16]), .B2(operand_1_x[17]), .B3(operand_1_x[16]), 
          .CI(mult_32u_32u_0_cin_lr_16), .CO(mco_120), .P0(mult_32u_32u_0_pp_8_17), 
          .P1(mult_32u_32u_0_pp_8_18)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_14_8 (.A0(muliplicand[16]), .A1(muliplicand[17]), 
          .A2(muliplicand[17]), .A3(muliplicand[18]), .B0(operand_1_x[15]), 
          .B1(operand_1_x[14]), .B2(operand_1_x[15]), .B3(operand_1_x[14]), 
          .CI(mco_112), .P0(mult_32u_32u_0_pp_7_31), .P1(mult_32u_32u_0_pp_7_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_14_7 (.A0(muliplicand[14]), .A1(muliplicand[15]), 
          .A2(muliplicand[15]), .A3(muliplicand[16]), .B0(operand_1_x[15]), 
          .B1(operand_1_x[14]), .B2(operand_1_x[15]), .B3(operand_1_x[14]), 
          .CI(mco_111), .CO(mco_112), .P0(mult_32u_32u_0_pp_7_29), .P1(mult_32u_32u_0_pp_7_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_14_6 (.A0(muliplicand[12]), .A1(muliplicand[13]), 
          .A2(muliplicand[13]), .A3(muliplicand[14]), .B0(operand_1_x[15]), 
          .B1(operand_1_x[14]), .B2(operand_1_x[15]), .B3(operand_1_x[14]), 
          .CI(mco_110), .CO(mco_111), .P0(mult_32u_32u_0_pp_7_27), .P1(mult_32u_32u_0_pp_7_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1S3AX result_i21 (.D(product[21]), .CK(w_clk_cpu), .Q(multiplier_result_w[21])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i21.GSR = "ENABLED";
    MULT2 mult_32u_32u_0_mult_14_5 (.A0(muliplicand[10]), .A1(muliplicand[11]), 
          .A2(muliplicand[11]), .A3(muliplicand[12]), .B0(operand_1_x[15]), 
          .B1(operand_1_x[14]), .B2(operand_1_x[15]), .B3(operand_1_x[14]), 
          .CI(mco_109), .CO(mco_110), .P0(mult_32u_32u_0_pp_7_25), .P1(mult_32u_32u_0_pp_7_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_14_4 (.A0(muliplicand[8]), .A1(muliplicand[9]), 
          .A2(muliplicand[9]), .A3(muliplicand[10]), .B0(operand_1_x[15]), 
          .B1(operand_1_x[14]), .B2(operand_1_x[15]), .B3(operand_1_x[14]), 
          .CI(mco_108), .CO(mco_109), .P0(mult_32u_32u_0_pp_7_23), .P1(mult_32u_32u_0_pp_7_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_14_3 (.A0(muliplicand[6]), .A1(muliplicand[7]), 
          .A2(muliplicand[7]), .A3(muliplicand[8]), .B0(operand_1_x[15]), 
          .B1(operand_1_x[14]), .B2(operand_1_x[15]), .B3(operand_1_x[14]), 
          .CI(mco_107), .CO(mco_108), .P0(mult_32u_32u_0_pp_7_21), .P1(mult_32u_32u_0_pp_7_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_14_2 (.A0(muliplicand[4]), .A1(muliplicand[5]), 
          .A2(muliplicand[5]), .A3(muliplicand[6]), .B0(operand_1_x[15]), 
          .B1(operand_1_x[14]), .B2(operand_1_x[15]), .B3(operand_1_x[14]), 
          .CI(mco_106), .CO(mco_107), .P0(mult_32u_32u_0_pp_7_19), .P1(mult_32u_32u_0_pp_7_20)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_14_1 (.A0(muliplicand[2]), .A1(muliplicand[3]), 
          .A2(muliplicand[3]), .A3(muliplicand[4]), .B0(operand_1_x[15]), 
          .B1(operand_1_x[14]), .B2(operand_1_x[15]), .B3(operand_1_x[14]), 
          .CI(mco_105), .CO(mco_106), .P0(mult_32u_32u_0_pp_7_17), .P1(mult_32u_32u_0_pp_7_18)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1S3AX result_i20 (.D(product[20]), .CK(w_clk_cpu), .Q(multiplier_result_w[20])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i20.GSR = "ENABLED";
    MULT2 mult_32u_32u_0_mult_14_0 (.A0(muliplicand[0]), .A1(muliplicand[1]), 
          .A2(muliplicand[1]), .A3(muliplicand[2]), .B0(operand_1_x[15]), 
          .B1(operand_1_x[14]), .B2(operand_1_x[15]), .B3(operand_1_x[14]), 
          .CI(mult_32u_32u_0_cin_lr_14), .CO(mco_105), .P0(mult_32u_32u_0_pp_7_15), 
          .P1(mult_32u_32u_0_pp_7_16)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_12_9 (.A0(muliplicand[18]), .A1(muliplicand[19]), 
          .A2(muliplicand[19]), .A3(muliplicand[20]), .B0(operand_1_x[13]), 
          .B1(operand_1_x[12]), .B2(operand_1_x[13]), .B3(operand_1_x[12]), 
          .CI(mco_98), .P0(mult_32u_32u_0_pp_6_31), .P1(mult_32u_32u_0_pp_6_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_12_8 (.A0(muliplicand[16]), .A1(muliplicand[17]), 
          .A2(muliplicand[17]), .A3(muliplicand[18]), .B0(operand_1_x[13]), 
          .B1(operand_1_x[12]), .B2(operand_1_x[13]), .B3(operand_1_x[12]), 
          .CI(mco_97), .CO(mco_98), .P0(mult_32u_32u_0_pp_6_29), .P1(mult_32u_32u_0_pp_6_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_12_7 (.A0(muliplicand[14]), .A1(muliplicand[15]), 
          .A2(muliplicand[15]), .A3(muliplicand[16]), .B0(operand_1_x[13]), 
          .B1(operand_1_x[12]), .B2(operand_1_x[13]), .B3(operand_1_x[12]), 
          .CI(mco_96), .CO(mco_97), .P0(mult_32u_32u_0_pp_6_27), .P1(mult_32u_32u_0_pp_6_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_12_6 (.A0(muliplicand[12]), .A1(muliplicand[13]), 
          .A2(muliplicand[13]), .A3(muliplicand[14]), .B0(operand_1_x[13]), 
          .B1(operand_1_x[12]), .B2(operand_1_x[13]), .B3(operand_1_x[12]), 
          .CI(mco_95), .CO(mco_96), .P0(mult_32u_32u_0_pp_6_25), .P1(mult_32u_32u_0_pp_6_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_12_5 (.A0(muliplicand[10]), .A1(muliplicand[11]), 
          .A2(muliplicand[11]), .A3(muliplicand[12]), .B0(operand_1_x[13]), 
          .B1(operand_1_x[12]), .B2(operand_1_x[13]), .B3(operand_1_x[12]), 
          .CI(mco_94), .CO(mco_95), .P0(mult_32u_32u_0_pp_6_23), .P1(mult_32u_32u_0_pp_6_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_12_4 (.A0(muliplicand[8]), .A1(muliplicand[9]), 
          .A2(muliplicand[9]), .A3(muliplicand[10]), .B0(operand_1_x[13]), 
          .B1(operand_1_x[12]), .B2(operand_1_x[13]), .B3(operand_1_x[12]), 
          .CI(mco_93), .CO(mco_94), .P0(mult_32u_32u_0_pp_6_21), .P1(mult_32u_32u_0_pp_6_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_12_3 (.A0(muliplicand[6]), .A1(muliplicand[7]), 
          .A2(muliplicand[7]), .A3(muliplicand[8]), .B0(operand_1_x[13]), 
          .B1(operand_1_x[12]), .B2(operand_1_x[13]), .B3(operand_1_x[12]), 
          .CI(mco_92), .CO(mco_93), .P0(mult_32u_32u_0_pp_6_19), .P1(mult_32u_32u_0_pp_6_20)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1S3AX result_i19 (.D(product[19]), .CK(w_clk_cpu), .Q(multiplier_result_w[19])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i19.GSR = "ENABLED";
    MULT2 mult_32u_32u_0_mult_12_2 (.A0(muliplicand[4]), .A1(muliplicand[5]), 
          .A2(muliplicand[5]), .A3(muliplicand[6]), .B0(operand_1_x[13]), 
          .B1(operand_1_x[12]), .B2(operand_1_x[13]), .B3(operand_1_x[12]), 
          .CI(mco_91), .CO(mco_92), .P0(mult_32u_32u_0_pp_6_17), .P1(mult_32u_32u_0_pp_6_18)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_12_1 (.A0(muliplicand[2]), .A1(muliplicand[3]), 
          .A2(muliplicand[3]), .A3(muliplicand[4]), .B0(operand_1_x[13]), 
          .B1(operand_1_x[12]), .B2(operand_1_x[13]), .B3(operand_1_x[12]), 
          .CI(mco_90), .CO(mco_91), .P0(mult_32u_32u_0_pp_6_15), .P1(mult_32u_32u_0_pp_6_16)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_12_0 (.A0(muliplicand[0]), .A1(muliplicand[1]), 
          .A2(muliplicand[1]), .A3(muliplicand[2]), .B0(operand_1_x[13]), 
          .B1(operand_1_x[12]), .B2(operand_1_x[13]), .B3(operand_1_x[12]), 
          .CI(mult_32u_32u_0_cin_lr_12), .CO(mco_90), .P0(mult_32u_32u_0_pp_6_13), 
          .P1(mult_32u_32u_0_pp_6_14)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1S3AX result_i18 (.D(product[18]), .CK(w_clk_cpu), .Q(multiplier_result_w[18])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i18.GSR = "ENABLED";
    MULT2 mult_32u_32u_0_mult_10_10 (.A0(muliplicand[20]), .A1(muliplicand[21]), 
          .A2(muliplicand[21]), .A3(muliplicand[22]), .B0(operand_1_x[11]), 
          .B1(operand_1_x[10]), .B2(operand_1_x[11]), .B3(operand_1_x[10]), 
          .CI(mco_84), .P0(mult_32u_32u_0_pp_5_31), .P1(mult_32u_32u_0_pp_5_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_10_9 (.A0(muliplicand[18]), .A1(muliplicand[19]), 
          .A2(muliplicand[19]), .A3(muliplicand[20]), .B0(operand_1_x[11]), 
          .B1(operand_1_x[10]), .B2(operand_1_x[11]), .B3(operand_1_x[10]), 
          .CI(mco_83), .CO(mco_84), .P0(mult_32u_32u_0_pp_5_29), .P1(mult_32u_32u_0_pp_5_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_10_8 (.A0(muliplicand[16]), .A1(muliplicand[17]), 
          .A2(muliplicand[17]), .A3(muliplicand[18]), .B0(operand_1_x[11]), 
          .B1(operand_1_x[10]), .B2(operand_1_x[11]), .B3(operand_1_x[10]), 
          .CI(mco_82), .CO(mco_83), .P0(mult_32u_32u_0_pp_5_27), .P1(mult_32u_32u_0_pp_5_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_10_7 (.A0(muliplicand[14]), .A1(muliplicand[15]), 
          .A2(muliplicand[15]), .A3(muliplicand[16]), .B0(operand_1_x[11]), 
          .B1(operand_1_x[10]), .B2(operand_1_x[11]), .B3(operand_1_x[10]), 
          .CI(mco_81), .CO(mco_82), .P0(mult_32u_32u_0_pp_5_25), .P1(mult_32u_32u_0_pp_5_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_10_6 (.A0(muliplicand[12]), .A1(muliplicand[13]), 
          .A2(muliplicand[13]), .A3(muliplicand[14]), .B0(operand_1_x[11]), 
          .B1(operand_1_x[10]), .B2(operand_1_x[11]), .B3(operand_1_x[10]), 
          .CI(mco_80), .CO(mco_81), .P0(mult_32u_32u_0_pp_5_23), .P1(mult_32u_32u_0_pp_5_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_10_5 (.A0(muliplicand[10]), .A1(muliplicand[11]), 
          .A2(muliplicand[11]), .A3(muliplicand[12]), .B0(operand_1_x[11]), 
          .B1(operand_1_x[10]), .B2(operand_1_x[11]), .B3(operand_1_x[10]), 
          .CI(mco_79), .CO(mco_80), .P0(mult_32u_32u_0_pp_5_21), .P1(mult_32u_32u_0_pp_5_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_10_4 (.A0(muliplicand[8]), .A1(muliplicand[9]), 
          .A2(muliplicand[9]), .A3(muliplicand[10]), .B0(operand_1_x[11]), 
          .B1(operand_1_x[10]), .B2(operand_1_x[11]), .B3(operand_1_x[10]), 
          .CI(mco_78), .CO(mco_79), .P0(mult_32u_32u_0_pp_5_19), .P1(mult_32u_32u_0_pp_5_20)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_10_3 (.A0(muliplicand[6]), .A1(muliplicand[7]), 
          .A2(muliplicand[7]), .A3(muliplicand[8]), .B0(operand_1_x[11]), 
          .B1(operand_1_x[10]), .B2(operand_1_x[11]), .B3(operand_1_x[10]), 
          .CI(mco_77), .CO(mco_78), .P0(mult_32u_32u_0_pp_5_17), .P1(mult_32u_32u_0_pp_5_18)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_10_2 (.A0(muliplicand[4]), .A1(muliplicand[5]), 
          .A2(muliplicand[5]), .A3(muliplicand[6]), .B0(operand_1_x[11]), 
          .B1(operand_1_x[10]), .B2(operand_1_x[11]), .B3(operand_1_x[10]), 
          .CI(mco_76), .CO(mco_77), .P0(mult_32u_32u_0_pp_5_15), .P1(mult_32u_32u_0_pp_5_16)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_10_1 (.A0(muliplicand[2]), .A1(muliplicand[3]), 
          .A2(muliplicand[3]), .A3(muliplicand[4]), .B0(operand_1_x[11]), 
          .B1(operand_1_x[10]), .B2(operand_1_x[11]), .B3(operand_1_x[10]), 
          .CI(mco_75), .CO(mco_76), .P0(mult_32u_32u_0_pp_5_13), .P1(mult_32u_32u_0_pp_5_14)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_10_0 (.A0(muliplicand[0]), .A1(muliplicand[1]), 
          .A2(muliplicand[1]), .A3(muliplicand[2]), .B0(operand_1_x[11]), 
          .B1(operand_1_x[10]), .B2(operand_1_x[11]), .B3(operand_1_x[10]), 
          .CI(mult_32u_32u_0_cin_lr_10), .CO(mco_75), .P0(mult_32u_32u_0_pp_5_11), 
          .P1(mult_32u_32u_0_pp_5_12)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B Cadd_mult_32u_32u_0_6_1 (.A0(GND_net), .A1(mult_32u_32u_0_pp_12_26), 
           .B0(GND_net), .B1(mult_32u_32u_0_pp_13_26), .CI(GND_net), .COUT(co_mult_32u_32u_0_6_1), 
           .S1(s_mult_32u_32u_0_6_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_8_11 (.A0(muliplicand[22]), .A1(muliplicand[23]), 
          .A2(muliplicand[23]), .A3(muliplicand[24]), .B0(operand_1_x[9]), 
          .B1(operand_1_x[8]), .B2(operand_1_x[9]), .B3(operand_1_x[8]), 
          .CI(mco_70), .P0(mult_32u_32u_0_pp_4_31), .P1(mult_32u_32u_0_pp_4_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_8_10 (.A0(muliplicand[20]), .A1(muliplicand[21]), 
          .A2(muliplicand[21]), .A3(muliplicand[22]), .B0(operand_1_x[9]), 
          .B1(operand_1_x[8]), .B2(operand_1_x[9]), .B3(operand_1_x[8]), 
          .CI(mco_69), .CO(mco_70), .P0(mult_32u_32u_0_pp_4_29), .P1(mult_32u_32u_0_pp_4_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_8_9 (.A0(muliplicand[18]), .A1(muliplicand[19]), 
          .A2(muliplicand[19]), .A3(muliplicand[20]), .B0(operand_1_x[9]), 
          .B1(operand_1_x[8]), .B2(operand_1_x[9]), .B3(operand_1_x[8]), 
          .CI(mco_68), .CO(mco_69), .P0(mult_32u_32u_0_pp_4_27), .P1(mult_32u_32u_0_pp_4_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_8_8 (.A0(muliplicand[16]), .A1(muliplicand[17]), 
          .A2(muliplicand[17]), .A3(muliplicand[18]), .B0(operand_1_x[9]), 
          .B1(operand_1_x[8]), .B2(operand_1_x[9]), .B3(operand_1_x[8]), 
          .CI(mco_67), .CO(mco_68), .P0(mult_32u_32u_0_pp_4_25), .P1(mult_32u_32u_0_pp_4_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_8_7 (.A0(muliplicand[14]), .A1(muliplicand[15]), 
          .A2(muliplicand[15]), .A3(muliplicand[16]), .B0(operand_1_x[9]), 
          .B1(operand_1_x[8]), .B2(operand_1_x[9]), .B3(operand_1_x[8]), 
          .CI(mco_66), .CO(mco_67), .P0(mult_32u_32u_0_pp_4_23), .P1(mult_32u_32u_0_pp_4_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_8_6 (.A0(muliplicand[12]), .A1(muliplicand[13]), 
          .A2(muliplicand[13]), .A3(muliplicand[14]), .B0(operand_1_x[9]), 
          .B1(operand_1_x[8]), .B2(operand_1_x[9]), .B3(operand_1_x[8]), 
          .CI(mco_65), .CO(mco_66), .P0(mult_32u_32u_0_pp_4_21), .P1(mult_32u_32u_0_pp_4_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_8_5 (.A0(muliplicand[10]), .A1(muliplicand[11]), 
          .A2(muliplicand[11]), .A3(muliplicand[12]), .B0(operand_1_x[9]), 
          .B1(operand_1_x[8]), .B2(operand_1_x[9]), .B3(operand_1_x[8]), 
          .CI(mco_64), .CO(mco_65), .P0(mult_32u_32u_0_pp_4_19), .P1(mult_32u_32u_0_pp_4_20)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_8_4 (.A0(muliplicand[8]), .A1(muliplicand[9]), 
          .A2(muliplicand[9]), .A3(muliplicand[10]), .B0(operand_1_x[9]), 
          .B1(operand_1_x[8]), .B2(operand_1_x[9]), .B3(operand_1_x[8]), 
          .CI(mco_63), .CO(mco_64), .P0(mult_32u_32u_0_pp_4_17), .P1(mult_32u_32u_0_pp_4_18)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_8_3 (.A0(muliplicand[6]), .A1(muliplicand[7]), 
          .A2(muliplicand[7]), .A3(muliplicand[8]), .B0(operand_1_x[9]), 
          .B1(operand_1_x[8]), .B2(operand_1_x[9]), .B3(operand_1_x[8]), 
          .CI(mco_62), .CO(mco_63), .P0(mult_32u_32u_0_pp_4_15), .P1(mult_32u_32u_0_pp_4_16)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_8_2 (.A0(muliplicand[4]), .A1(muliplicand[5]), 
          .A2(muliplicand[5]), .A3(muliplicand[6]), .B0(operand_1_x[9]), 
          .B1(operand_1_x[8]), .B2(operand_1_x[9]), .B3(operand_1_x[8]), 
          .CI(mco_61), .CO(mco_62), .P0(mult_32u_32u_0_pp_4_13), .P1(mult_32u_32u_0_pp_4_14)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_8_1 (.A0(muliplicand[2]), .A1(muliplicand[3]), 
          .A2(muliplicand[3]), .A3(muliplicand[4]), .B0(operand_1_x[9]), 
          .B1(operand_1_x[8]), .B2(operand_1_x[9]), .B3(operand_1_x[8]), 
          .CI(mco_60), .CO(mco_61), .P0(mult_32u_32u_0_pp_4_11), .P1(mult_32u_32u_0_pp_4_12)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_8_0 (.A0(muliplicand[0]), .A1(muliplicand[1]), 
          .A2(muliplicand[1]), .A3(muliplicand[2]), .B0(operand_1_x[9]), 
          .B1(operand_1_x[8]), .B2(operand_1_x[9]), .B3(operand_1_x[8]), 
          .CI(mult_32u_32u_0_cin_lr_8), .CO(mco_60), .P0(mult_32u_32u_0_pp_4_9), 
          .P1(mult_32u_32u_0_pp_4_10)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1S3AX result_i17 (.D(product[17]), .CK(w_clk_cpu), .Q(multiplier_result_w[17])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i17.GSR = "ENABLED";
    MULT2 mult_32u_32u_0_mult_6_12 (.A0(muliplicand[24]), .A1(muliplicand[25]), 
          .A2(muliplicand[25]), .A3(muliplicand[26]), .B0(operand_1_x[7]), 
          .B1(operand_1_x[6]), .B2(operand_1_x[7]), .B3(operand_1_x[6]), 
          .CI(mco_56), .P0(mult_32u_32u_0_pp_3_31), .P1(mult_32u_32u_0_pp_3_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_6_11 (.A0(muliplicand[22]), .A1(muliplicand[23]), 
          .A2(muliplicand[23]), .A3(muliplicand[24]), .B0(operand_1_x[7]), 
          .B1(operand_1_x[6]), .B2(operand_1_x[7]), .B3(operand_1_x[6]), 
          .CI(mco_55), .CO(mco_56), .P0(mult_32u_32u_0_pp_3_29), .P1(mult_32u_32u_0_pp_3_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_6_10 (.A0(muliplicand[20]), .A1(muliplicand[21]), 
          .A2(muliplicand[21]), .A3(muliplicand[22]), .B0(operand_1_x[7]), 
          .B1(operand_1_x[6]), .B2(operand_1_x[7]), .B3(operand_1_x[6]), 
          .CI(mco_54), .CO(mco_55), .P0(mult_32u_32u_0_pp_3_27), .P1(mult_32u_32u_0_pp_3_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_6_9 (.A0(muliplicand[18]), .A1(muliplicand[19]), 
          .A2(muliplicand[19]), .A3(muliplicand[20]), .B0(operand_1_x[7]), 
          .B1(operand_1_x[6]), .B2(operand_1_x[7]), .B3(operand_1_x[6]), 
          .CI(mco_53), .CO(mco_54), .P0(mult_32u_32u_0_pp_3_25), .P1(mult_32u_32u_0_pp_3_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_6_8 (.A0(muliplicand[16]), .A1(muliplicand[17]), 
          .A2(muliplicand[17]), .A3(muliplicand[18]), .B0(operand_1_x[7]), 
          .B1(operand_1_x[6]), .B2(operand_1_x[7]), .B3(operand_1_x[6]), 
          .CI(mco_52), .CO(mco_53), .P0(mult_32u_32u_0_pp_3_23), .P1(mult_32u_32u_0_pp_3_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_6_7 (.A0(muliplicand[14]), .A1(muliplicand[15]), 
          .A2(muliplicand[15]), .A3(muliplicand[16]), .B0(operand_1_x[7]), 
          .B1(operand_1_x[6]), .B2(operand_1_x[7]), .B3(operand_1_x[6]), 
          .CI(mco_51), .CO(mco_52), .P0(mult_32u_32u_0_pp_3_21), .P1(mult_32u_32u_0_pp_3_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_6_6 (.A0(muliplicand[12]), .A1(muliplicand[13]), 
          .A2(muliplicand[13]), .A3(muliplicand[14]), .B0(operand_1_x[7]), 
          .B1(operand_1_x[6]), .B2(operand_1_x[7]), .B3(operand_1_x[6]), 
          .CI(mco_50), .CO(mco_51), .P0(mult_32u_32u_0_pp_3_19), .P1(mult_32u_32u_0_pp_3_20)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_6_5 (.A0(muliplicand[10]), .A1(muliplicand[11]), 
          .A2(muliplicand[11]), .A3(muliplicand[12]), .B0(operand_1_x[7]), 
          .B1(operand_1_x[6]), .B2(operand_1_x[7]), .B3(operand_1_x[6]), 
          .CI(mco_49), .CO(mco_50), .P0(mult_32u_32u_0_pp_3_17), .P1(mult_32u_32u_0_pp_3_18)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_6_4 (.A0(muliplicand[8]), .A1(muliplicand[9]), 
          .A2(muliplicand[9]), .A3(muliplicand[10]), .B0(operand_1_x[7]), 
          .B1(operand_1_x[6]), .B2(operand_1_x[7]), .B3(operand_1_x[6]), 
          .CI(mco_48), .CO(mco_49), .P0(mult_32u_32u_0_pp_3_15), .P1(mult_32u_32u_0_pp_3_16)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_6_3 (.A0(muliplicand[6]), .A1(muliplicand[7]), 
          .A2(muliplicand[7]), .A3(muliplicand[8]), .B0(operand_1_x[7]), 
          .B1(operand_1_x[6]), .B2(operand_1_x[7]), .B3(operand_1_x[6]), 
          .CI(mco_47), .CO(mco_48), .P0(mult_32u_32u_0_pp_3_13), .P1(mult_32u_32u_0_pp_3_14)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_6_2 (.A0(muliplicand[4]), .A1(muliplicand[5]), 
          .A2(muliplicand[5]), .A3(muliplicand[6]), .B0(operand_1_x[7]), 
          .B1(operand_1_x[6]), .B2(operand_1_x[7]), .B3(operand_1_x[6]), 
          .CI(mco_46), .CO(mco_47), .P0(mult_32u_32u_0_pp_3_11), .P1(mult_32u_32u_0_pp_3_12)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_6_1 (.A0(muliplicand[2]), .A1(muliplicand[3]), 
          .A2(muliplicand[3]), .A3(muliplicand[4]), .B0(operand_1_x[7]), 
          .B1(operand_1_x[6]), .B2(operand_1_x[7]), .B3(operand_1_x[6]), 
          .CI(mco_45), .CO(mco_46), .P0(mult_32u_32u_0_pp_3_9), .P1(mult_32u_32u_0_pp_3_10)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_6_0 (.A0(muliplicand[0]), .A1(muliplicand[1]), 
          .A2(muliplicand[1]), .A3(muliplicand[2]), .B0(operand_1_x[7]), 
          .B1(operand_1_x[6]), .B2(operand_1_x[7]), .B3(operand_1_x[6]), 
          .CI(mult_32u_32u_0_cin_lr_6), .CO(mco_45), .P0(mult_32u_32u_0_pp_3_7), 
          .P1(mult_32u_32u_0_pp_3_8)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_4_13 (.A0(muliplicand[26]), .A1(muliplicand[27]), 
          .A2(muliplicand[27]), .A3(muliplicand[28]), .B0(operand_1_x[5]), 
          .B1(operand_1_x[4]), .B2(operand_1_x[5]), .B3(operand_1_x[4]), 
          .CI(mco_42), .P0(mult_32u_32u_0_pp_2_31), .P1(mult_32u_32u_0_pp_2_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_4_12 (.A0(muliplicand[24]), .A1(muliplicand[25]), 
          .A2(muliplicand[25]), .A3(muliplicand[26]), .B0(operand_1_x[5]), 
          .B1(operand_1_x[4]), .B2(operand_1_x[5]), .B3(operand_1_x[4]), 
          .CI(mco_41), .CO(mco_42), .P0(mult_32u_32u_0_pp_2_29), .P1(mult_32u_32u_0_pp_2_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1S3AX result_i16 (.D(product[16]), .CK(w_clk_cpu), .Q(multiplier_result_w[16])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i16.GSR = "ENABLED";
    MULT2 mult_32u_32u_0_mult_4_11 (.A0(muliplicand[22]), .A1(muliplicand[23]), 
          .A2(muliplicand[23]), .A3(muliplicand[24]), .B0(operand_1_x[5]), 
          .B1(operand_1_x[4]), .B2(operand_1_x[5]), .B3(operand_1_x[4]), 
          .CI(mco_40), .CO(mco_41), .P0(mult_32u_32u_0_pp_2_27), .P1(mult_32u_32u_0_pp_2_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_4_10 (.A0(muliplicand[20]), .A1(muliplicand[21]), 
          .A2(muliplicand[21]), .A3(muliplicand[22]), .B0(operand_1_x[5]), 
          .B1(operand_1_x[4]), .B2(operand_1_x[5]), .B3(operand_1_x[4]), 
          .CI(mco_39), .CO(mco_40), .P0(mult_32u_32u_0_pp_2_25), .P1(mult_32u_32u_0_pp_2_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_4_9 (.A0(muliplicand[18]), .A1(muliplicand[19]), 
          .A2(muliplicand[19]), .A3(muliplicand[20]), .B0(operand_1_x[5]), 
          .B1(operand_1_x[4]), .B2(operand_1_x[5]), .B3(operand_1_x[4]), 
          .CI(mco_38), .CO(mco_39), .P0(mult_32u_32u_0_pp_2_23), .P1(mult_32u_32u_0_pp_2_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_4_8 (.A0(muliplicand[16]), .A1(muliplicand[17]), 
          .A2(muliplicand[17]), .A3(muliplicand[18]), .B0(operand_1_x[5]), 
          .B1(operand_1_x[4]), .B2(operand_1_x[5]), .B3(operand_1_x[4]), 
          .CI(mco_37), .CO(mco_38), .P0(mult_32u_32u_0_pp_2_21), .P1(mult_32u_32u_0_pp_2_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_4_7 (.A0(muliplicand[14]), .A1(muliplicand[15]), 
          .A2(muliplicand[15]), .A3(muliplicand[16]), .B0(operand_1_x[5]), 
          .B1(operand_1_x[4]), .B2(operand_1_x[5]), .B3(operand_1_x[4]), 
          .CI(mco_36), .CO(mco_37), .P0(mult_32u_32u_0_pp_2_19), .P1(mult_32u_32u_0_pp_2_20)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_4_6 (.A0(muliplicand[12]), .A1(muliplicand[13]), 
          .A2(muliplicand[13]), .A3(muliplicand[14]), .B0(operand_1_x[5]), 
          .B1(operand_1_x[4]), .B2(operand_1_x[5]), .B3(operand_1_x[4]), 
          .CI(mco_35), .CO(mco_36), .P0(mult_32u_32u_0_pp_2_17), .P1(mult_32u_32u_0_pp_2_18)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_4_5 (.A0(muliplicand[10]), .A1(muliplicand[11]), 
          .A2(muliplicand[11]), .A3(muliplicand[12]), .B0(operand_1_x[5]), 
          .B1(operand_1_x[4]), .B2(operand_1_x[5]), .B3(operand_1_x[4]), 
          .CI(mco_34), .CO(mco_35), .P0(mult_32u_32u_0_pp_2_15), .P1(mult_32u_32u_0_pp_2_16)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_4_4 (.A0(muliplicand[8]), .A1(muliplicand[9]), 
          .A2(muliplicand[9]), .A3(muliplicand[10]), .B0(operand_1_x[5]), 
          .B1(operand_1_x[4]), .B2(operand_1_x[5]), .B3(operand_1_x[4]), 
          .CI(mco_33), .CO(mco_34), .P0(mult_32u_32u_0_pp_2_13), .P1(mult_32u_32u_0_pp_2_14)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_4_3 (.A0(muliplicand[6]), .A1(muliplicand[7]), 
          .A2(muliplicand[7]), .A3(muliplicand[8]), .B0(operand_1_x[5]), 
          .B1(operand_1_x[4]), .B2(operand_1_x[5]), .B3(operand_1_x[4]), 
          .CI(mco_32), .CO(mco_33), .P0(mult_32u_32u_0_pp_2_11), .P1(mult_32u_32u_0_pp_2_12)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_4_2 (.A0(muliplicand[4]), .A1(muliplicand[5]), 
          .A2(muliplicand[5]), .A3(muliplicand[6]), .B0(operand_1_x[5]), 
          .B1(operand_1_x[4]), .B2(operand_1_x[5]), .B3(operand_1_x[4]), 
          .CI(mco_31), .CO(mco_32), .P0(mult_32u_32u_0_pp_2_9), .P1(mult_32u_32u_0_pp_2_10)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_4_1 (.A0(muliplicand[2]), .A1(muliplicand[3]), 
          .A2(muliplicand[3]), .A3(muliplicand[4]), .B0(operand_1_x[5]), 
          .B1(operand_1_x[4]), .B2(operand_1_x[5]), .B3(operand_1_x[4]), 
          .CI(mco_30), .CO(mco_31), .P0(mult_32u_32u_0_pp_2_7), .P1(mult_32u_32u_0_pp_2_8)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_4_0 (.A0(muliplicand[0]), .A1(muliplicand[1]), 
          .A2(muliplicand[1]), .A3(muliplicand[2]), .B0(operand_1_x[5]), 
          .B1(operand_1_x[4]), .B2(operand_1_x[5]), .B3(operand_1_x[4]), 
          .CI(mult_32u_32u_0_cin_lr_4), .CO(mco_30), .P0(mult_32u_32u_0_pp_2_5), 
          .P1(mult_32u_32u_0_pp_2_6)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_2_14 (.A0(muliplicand[28]), .A1(muliplicand[29]), 
          .A2(muliplicand[29]), .A3(muliplicand[30]), .B0(operand_1_x[3]), 
          .B1(operand_1_x[2]), .B2(operand_1_x[3]), .B3(operand_1_x[2]), 
          .CI(mco_28), .P0(mult_32u_32u_0_pp_1_31), .P1(mult_32u_32u_0_pp_1_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_2_13 (.A0(muliplicand[26]), .A1(muliplicand[27]), 
          .A2(muliplicand[27]), .A3(muliplicand[28]), .B0(operand_1_x[3]), 
          .B1(operand_1_x[2]), .B2(operand_1_x[3]), .B3(operand_1_x[2]), 
          .CI(mco_27), .CO(mco_28), .P0(mult_32u_32u_0_pp_1_29), .P1(mult_32u_32u_0_pp_1_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_2_12 (.A0(muliplicand[24]), .A1(muliplicand[25]), 
          .A2(muliplicand[25]), .A3(muliplicand[26]), .B0(operand_1_x[3]), 
          .B1(operand_1_x[2]), .B2(operand_1_x[3]), .B3(operand_1_x[2]), 
          .CI(mco_26), .CO(mco_27), .P0(mult_32u_32u_0_pp_1_27), .P1(mult_32u_32u_0_pp_1_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1S3AX result_i15 (.D(product[15]), .CK(w_clk_cpu), .Q(multiplier_result_w[15])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i15.GSR = "ENABLED";
    MULT2 mult_32u_32u_0_mult_2_11 (.A0(muliplicand[22]), .A1(muliplicand[23]), 
          .A2(muliplicand[23]), .A3(muliplicand[24]), .B0(operand_1_x[3]), 
          .B1(operand_1_x[2]), .B2(operand_1_x[3]), .B3(operand_1_x[2]), 
          .CI(mco_25), .CO(mco_26), .P0(mult_32u_32u_0_pp_1_25), .P1(mult_32u_32u_0_pp_1_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_2_10 (.A0(muliplicand[20]), .A1(muliplicand[21]), 
          .A2(muliplicand[21]), .A3(muliplicand[22]), .B0(operand_1_x[3]), 
          .B1(operand_1_x[2]), .B2(operand_1_x[3]), .B3(operand_1_x[2]), 
          .CI(mco_24), .CO(mco_25), .P0(mult_32u_32u_0_pp_1_23), .P1(mult_32u_32u_0_pp_1_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_2_9 (.A0(muliplicand[18]), .A1(muliplicand[19]), 
          .A2(muliplicand[19]), .A3(muliplicand[20]), .B0(operand_1_x[3]), 
          .B1(operand_1_x[2]), .B2(operand_1_x[3]), .B3(operand_1_x[2]), 
          .CI(mco_23), .CO(mco_24), .P0(mult_32u_32u_0_pp_1_21), .P1(mult_32u_32u_0_pp_1_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_2_8 (.A0(muliplicand[16]), .A1(muliplicand[17]), 
          .A2(muliplicand[17]), .A3(muliplicand[18]), .B0(operand_1_x[3]), 
          .B1(operand_1_x[2]), .B2(operand_1_x[3]), .B3(operand_1_x[2]), 
          .CI(mco_22), .CO(mco_23), .P0(mult_32u_32u_0_pp_1_19), .P1(mult_32u_32u_0_pp_1_20)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_2_7 (.A0(muliplicand[14]), .A1(muliplicand[15]), 
          .A2(muliplicand[15]), .A3(muliplicand[16]), .B0(operand_1_x[3]), 
          .B1(operand_1_x[2]), .B2(operand_1_x[3]), .B3(operand_1_x[2]), 
          .CI(mco_21), .CO(mco_22), .P0(mult_32u_32u_0_pp_1_17), .P1(mult_32u_32u_0_pp_1_18)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_2_6 (.A0(muliplicand[12]), .A1(muliplicand[13]), 
          .A2(muliplicand[13]), .A3(muliplicand[14]), .B0(operand_1_x[3]), 
          .B1(operand_1_x[2]), .B2(operand_1_x[3]), .B3(operand_1_x[2]), 
          .CI(mco_20), .CO(mco_21), .P0(mult_32u_32u_0_pp_1_15), .P1(mult_32u_32u_0_pp_1_16)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_2_5 (.A0(muliplicand[10]), .A1(muliplicand[11]), 
          .A2(muliplicand[11]), .A3(muliplicand[12]), .B0(operand_1_x[3]), 
          .B1(operand_1_x[2]), .B2(operand_1_x[3]), .B3(operand_1_x[2]), 
          .CI(mco_19), .CO(mco_20), .P0(mult_32u_32u_0_pp_1_13), .P1(mult_32u_32u_0_pp_1_14)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_2_4 (.A0(muliplicand[8]), .A1(muliplicand[9]), 
          .A2(muliplicand[9]), .A3(muliplicand[10]), .B0(operand_1_x[3]), 
          .B1(operand_1_x[2]), .B2(operand_1_x[3]), .B3(operand_1_x[2]), 
          .CI(mco_18), .CO(mco_19), .P0(mult_32u_32u_0_pp_1_11), .P1(mult_32u_32u_0_pp_1_12)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_2_3 (.A0(muliplicand[6]), .A1(muliplicand[7]), 
          .A2(muliplicand[7]), .A3(muliplicand[8]), .B0(operand_1_x[3]), 
          .B1(operand_1_x[2]), .B2(operand_1_x[3]), .B3(operand_1_x[2]), 
          .CI(mco_17), .CO(mco_18), .P0(mult_32u_32u_0_pp_1_9), .P1(mult_32u_32u_0_pp_1_10)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_2_2 (.A0(muliplicand[4]), .A1(muliplicand[5]), 
          .A2(muliplicand[5]), .A3(muliplicand[6]), .B0(operand_1_x[3]), 
          .B1(operand_1_x[2]), .B2(operand_1_x[3]), .B3(operand_1_x[2]), 
          .CI(mco_16), .CO(mco_17), .P0(mult_32u_32u_0_pp_1_7), .P1(mult_32u_32u_0_pp_1_8)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_2_1 (.A0(muliplicand[2]), .A1(muliplicand[3]), 
          .A2(muliplicand[3]), .A3(muliplicand[4]), .B0(operand_1_x[3]), 
          .B1(operand_1_x[2]), .B2(operand_1_x[3]), .B3(operand_1_x[2]), 
          .CI(mco_15), .CO(mco_16), .P0(mult_32u_32u_0_pp_1_5), .P1(mult_32u_32u_0_pp_1_6)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_4_8 (.A0(mult_32u_32u_0_pp_8_31), .A1(mult_32u_32u_0_pp_8_32), 
           .B0(mult_32u_32u_0_pp_9_31), .B1(mult_32u_32u_0_pp_9_32), .CI(co_mult_32u_32u_0_4_7), 
           .S0(s_mult_32u_32u_0_4_31), .S1(s_mult_32u_32u_0_4_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_2_0 (.A0(muliplicand[0]), .A1(muliplicand[1]), 
          .A2(muliplicand[1]), .A3(muliplicand[2]), .B0(operand_1_x[3]), 
          .B1(operand_1_x[2]), .B2(operand_1_x[3]), .B3(operand_1_x[2]), 
          .CI(mult_32u_32u_0_cin_lr_2), .CO(mco_15), .P0(mult_32u_32u_0_pp_1_3), 
          .P1(mult_32u_32u_0_pp_1_4)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_0_15 (.A0(muliplicand[30]), .A1(muliplicand[31]), 
          .A2(muliplicand[31]), .A3(GND_net), .B0(operand_1_x[1]), .B1(operand_1_x[0]), 
          .B2(operand_1_x[1]), .B3(operand_1_x[0]), .CI(mco_14), .P0(mult_32u_32u_0_pp_0_31), 
          .P1(mult_32u_32u_0_pp_0_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_12_13 (.A0(s_mult_32u_32u_0_8_31), .A1(s_mult_32u_32u_0_8_32), 
           .B0(s_mult_32u_32u_0_9_31), .B1(s_mult_32u_32u_0_9_32), .CI(co_mult_32u_32u_0_12_12), 
           .S0(s_mult_32u_32u_0_12_31), .S1(s_mult_32u_32u_0_12_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_0_14 (.A0(muliplicand[28]), .A1(muliplicand[29]), 
          .A2(muliplicand[29]), .A3(muliplicand[30]), .B0(operand_1_x[1]), 
          .B1(operand_1_x[0]), .B2(operand_1_x[1]), .B3(operand_1_x[0]), 
          .CI(mco_13), .CO(mco_14), .P0(mult_32u_32u_0_pp_0_29), .P1(mult_32u_32u_0_pp_0_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_0_13 (.A0(muliplicand[26]), .A1(muliplicand[27]), 
          .A2(muliplicand[27]), .A3(muliplicand[28]), .B0(operand_1_x[1]), 
          .B1(operand_1_x[0]), .B2(operand_1_x[1]), .B3(operand_1_x[0]), 
          .CI(mco_12), .CO(mco_13), .P0(mult_32u_32u_0_pp_0_27), .P1(mult_32u_32u_0_pp_0_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_12_12 (.A0(s_mult_32u_32u_0_8_29), .A1(s_mult_32u_32u_0_8_30), 
           .B0(s_mult_32u_32u_0_9_29), .B1(s_mult_32u_32u_0_9_30), .CI(co_mult_32u_32u_0_12_11), 
           .COUT(co_mult_32u_32u_0_12_12), .S0(s_mult_32u_32u_0_12_29), 
           .S1(s_mult_32u_32u_0_12_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_12_11 (.A0(s_mult_32u_32u_0_8_27), .A1(s_mult_32u_32u_0_8_28), 
           .B0(s_mult_32u_32u_0_9_27), .B1(s_mult_32u_32u_0_9_28), .CI(co_mult_32u_32u_0_12_10), 
           .COUT(co_mult_32u_32u_0_12_11), .S0(s_mult_32u_32u_0_12_27), 
           .S1(s_mult_32u_32u_0_12_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_4_7 (.A0(mult_32u_32u_0_pp_8_29), .A1(mult_32u_32u_0_pp_8_30), 
           .B0(mult_32u_32u_0_pp_9_29), .B1(mult_32u_32u_0_pp_9_30), .CI(co_mult_32u_32u_0_4_6), 
           .COUT(co_mult_32u_32u_0_4_7), .S0(s_mult_32u_32u_0_4_29), .S1(s_mult_32u_32u_0_4_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B Cadd_mult_32u_32u_0_5_1 (.A0(GND_net), .A1(mult_32u_32u_0_pp_10_22), 
           .B0(GND_net), .B1(mult_32u_32u_0_pp_11_22), .CI(GND_net), .COUT(co_mult_32u_32u_0_5_1), 
           .S1(s_mult_32u_32u_0_5_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_0_12 (.A0(muliplicand[24]), .A1(muliplicand[25]), 
          .A2(muliplicand[25]), .A3(muliplicand[26]), .B0(operand_1_x[1]), 
          .B1(operand_1_x[0]), .B2(operand_1_x[1]), .B3(operand_1_x[0]), 
          .CI(mco_11), .CO(mco_12), .P0(mult_32u_32u_0_pp_0_25), .P1(mult_32u_32u_0_pp_0_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_12_10 (.A0(s_mult_32u_32u_0_8_25), .A1(s_mult_32u_32u_0_8_26), 
           .B0(s_mult_32u_32u_0_9_25), .B1(s_mult_32u_32u_0_9_26), .CI(co_mult_32u_32u_0_12_9), 
           .COUT(co_mult_32u_32u_0_12_10), .S0(s_mult_32u_32u_0_12_25), 
           .S1(s_mult_32u_32u_0_12_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_12_9 (.A0(s_mult_32u_32u_0_8_23), .A1(s_mult_32u_32u_0_8_24), 
           .B0(s_mult_32u_32u_0_9_23), .B1(s_mult_32u_32u_0_9_24), .CI(co_mult_32u_32u_0_12_8), 
           .COUT(co_mult_32u_32u_0_12_9), .S0(s_mult_32u_32u_0_12_23), .S1(s_mult_32u_32u_0_12_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_4_6 (.A0(mult_32u_32u_0_pp_8_27), .A1(mult_32u_32u_0_pp_8_28), 
           .B0(mult_32u_32u_0_pp_9_27), .B1(mult_32u_32u_0_pp_9_28), .CI(co_mult_32u_32u_0_4_5), 
           .COUT(co_mult_32u_32u_0_4_6), .S0(s_mult_32u_32u_0_4_27), .S1(s_mult_32u_32u_0_4_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_4_5 (.A0(mult_32u_32u_0_pp_8_25), .A1(mult_32u_32u_0_pp_8_26), 
           .B0(mult_32u_32u_0_pp_9_25), .B1(mult_32u_32u_0_pp_9_26), .CI(co_mult_32u_32u_0_4_4), 
           .COUT(co_mult_32u_32u_0_4_5), .S0(s_mult_32u_32u_0_4_25), .S1(s_mult_32u_32u_0_4_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_12_8 (.A0(s_mult_32u_32u_0_8_21), .A1(s_mult_32u_32u_0_8_22), 
           .B0(s_mult_32u_32u_0_9_21), .B1(s_mult_32u_32u_0_9_22), .CI(co_mult_32u_32u_0_12_7), 
           .COUT(co_mult_32u_32u_0_12_8), .S0(s_mult_32u_32u_0_12_21), .S1(s_mult_32u_32u_0_12_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_4_4 (.A0(mult_32u_32u_0_pp_8_23), .A1(mult_32u_32u_0_pp_8_24), 
           .B0(mult_32u_32u_0_pp_9_23), .B1(mult_32u_32u_0_pp_9_24), .CI(co_mult_32u_32u_0_4_3), 
           .COUT(co_mult_32u_32u_0_4_4), .S0(s_mult_32u_32u_0_4_23), .S1(s_mult_32u_32u_0_4_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_4_3 (.A0(mult_32u_32u_0_pp_8_21), .A1(mult_32u_32u_0_pp_8_22), 
           .B0(mult_32u_32u_0_pp_9_21), .B1(mult_32u_32u_0_pp_9_22), .CI(co_mult_32u_32u_0_4_2), 
           .COUT(co_mult_32u_32u_0_4_3), .S0(s_mult_32u_32u_0_4_21), .S1(s_mult_32u_32u_0_4_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_4_2 (.A0(mult_32u_32u_0_pp_8_19), .A1(mult_32u_32u_0_pp_8_20), 
           .B0(mult_32u_32u_0_pp_9_19), .B1(mult_32u_32u_0_pp_9_20), .CI(co_mult_32u_32u_0_4_1), 
           .COUT(co_mult_32u_32u_0_4_2), .S0(s_mult_32u_32u_0_4_19), .S1(s_mult_32u_32u_0_4_20)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_12_7 (.A0(s_mult_32u_32u_0_8_19), .A1(s_mult_32u_32u_0_8_20), 
           .B0(s_mult_32u_32u_0_9_19), .B1(s_mult_32u_32u_0_9_20), .CI(co_mult_32u_32u_0_12_6), 
           .COUT(co_mult_32u_32u_0_12_7), .S0(s_mult_32u_32u_0_12_19), .S1(s_mult_32u_32u_0_12_20)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_12_6 (.A0(s_mult_32u_32u_0_8_17), .A1(s_mult_32u_32u_0_8_18), 
           .B0(s_mult_32u_32u_0_9_17), .B1(s_mult_32u_32u_0_9_18), .CI(co_mult_32u_32u_0_12_5), 
           .COUT(co_mult_32u_32u_0_12_6), .S0(s_mult_32u_32u_0_12_17), .S1(s_mult_32u_32u_0_12_18)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B Cadd_mult_32u_32u_0_4_1 (.A0(GND_net), .A1(mult_32u_32u_0_pp_8_18), 
           .B0(GND_net), .B1(mult_32u_32u_0_pp_9_18), .CI(GND_net), .COUT(co_mult_32u_32u_0_4_1), 
           .S1(s_mult_32u_32u_0_4_18)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_0_11 (.A0(muliplicand[22]), .A1(muliplicand[23]), 
          .A2(muliplicand[23]), .A3(muliplicand[24]), .B0(operand_1_x[1]), 
          .B1(operand_1_x[0]), .B2(operand_1_x[1]), .B3(operand_1_x[0]), 
          .CI(mco_10), .CO(mco_11), .P0(mult_32u_32u_0_pp_0_23), .P1(mult_32u_32u_0_pp_0_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_12_5 (.A0(s_mult_32u_32u_0_8_15), .A1(s_mult_32u_32u_0_8_16), 
           .B0(s_mult_32u_32u_0_9_15), .B1(s_mult_32u_32u_0_9_16), .CI(co_mult_32u_32u_0_12_4), 
           .COUT(co_mult_32u_32u_0_12_5), .S0(product_31__N_2324[15]), .S1(s_mult_32u_32u_0_12_16)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_0_10 (.A0(muliplicand[20]), .A1(muliplicand[21]), 
          .A2(muliplicand[21]), .A3(muliplicand[22]), .B0(operand_1_x[1]), 
          .B1(operand_1_x[0]), .B2(operand_1_x[1]), .B3(operand_1_x[0]), 
          .CI(mco_9), .CO(mco_10), .P0(mult_32u_32u_0_pp_0_21), .P1(mult_32u_32u_0_pp_0_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_0_9 (.A0(muliplicand[18]), .A1(muliplicand[19]), 
          .A2(muliplicand[19]), .A3(muliplicand[20]), .B0(operand_1_x[1]), 
          .B1(operand_1_x[0]), .B2(operand_1_x[1]), .B3(operand_1_x[0]), 
          .CI(mco_8), .CO(mco_9), .P0(mult_32u_32u_0_pp_0_19), .P1(mult_32u_32u_0_pp_0_20)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_0_8 (.A0(muliplicand[16]), .A1(muliplicand[17]), 
          .A2(muliplicand[17]), .A3(muliplicand[18]), .B0(operand_1_x[1]), 
          .B1(operand_1_x[0]), .B2(operand_1_x[1]), .B3(operand_1_x[0]), 
          .CI(mco_7), .CO(mco_8), .P0(mult_32u_32u_0_pp_0_17), .P1(mult_32u_32u_0_pp_0_18)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_0_7 (.A0(muliplicand[14]), .A1(muliplicand[15]), 
          .A2(muliplicand[15]), .A3(muliplicand[16]), .B0(operand_1_x[1]), 
          .B1(operand_1_x[0]), .B2(operand_1_x[1]), .B3(operand_1_x[0]), 
          .CI(mco_6), .CO(mco_7), .P0(mult_32u_32u_0_pp_0_15), .P1(mult_32u_32u_0_pp_0_16)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_0_6 (.A0(muliplicand[12]), .A1(muliplicand[13]), 
          .A2(muliplicand[13]), .A3(muliplicand[14]), .B0(operand_1_x[1]), 
          .B1(operand_1_x[0]), .B2(operand_1_x[1]), .B3(operand_1_x[0]), 
          .CI(mco_5), .CO(mco_6), .P0(mult_32u_32u_0_pp_0_13), .P1(mult_32u_32u_0_pp_0_14)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_12_4 (.A0(s_mult_32u_32u_0_8_13), .A1(s_mult_32u_32u_0_8_14), 
           .B0(s_mult_32u_32u_0_9_13), .B1(s_mult_32u_32u_0_9_14), .CI(co_mult_32u_32u_0_12_3), 
           .COUT(co_mult_32u_32u_0_12_4), .S0(product_31__N_2324[13]), .S1(product_31__N_2324[14])) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_0_5 (.A0(muliplicand[10]), .A1(muliplicand[11]), 
          .A2(muliplicand[11]), .A3(muliplicand[12]), .B0(operand_1_x[1]), 
          .B1(operand_1_x[0]), .B2(operand_1_x[1]), .B3(operand_1_x[0]), 
          .CI(mco_4), .CO(mco_5), .P0(mult_32u_32u_0_pp_0_11), .P1(mult_32u_32u_0_pp_0_12)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_12_3 (.A0(s_mult_32u_32u_0_8_11), .A1(s_mult_32u_32u_0_8_12), 
           .B0(s_mult_32u_32u_0_2_11), .B1(s_mult_32u_32u_0_9_12), .CI(co_mult_32u_32u_0_12_2), 
           .COUT(co_mult_32u_32u_0_12_3), .S0(product_31__N_2324[11]), .S1(product_31__N_2324[12])) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_0_4 (.A0(muliplicand[8]), .A1(muliplicand[9]), 
          .A2(muliplicand[9]), .A3(muliplicand[10]), .B0(operand_1_x[1]), 
          .B1(operand_1_x[0]), .B2(operand_1_x[1]), .B3(operand_1_x[0]), 
          .CI(mco_3), .CO(mco_4), .P0(mult_32u_32u_0_pp_0_9), .P1(mult_32u_32u_0_pp_0_10)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_12_2 (.A0(s_mult_32u_32u_0_8_9), .A1(s_mult_32u_32u_0_8_10), 
           .B0(mult_32u_32u_0_pp_4_9), .B1(s_mult_32u_32u_0_2_10), .CI(co_mult_32u_32u_0_12_1), 
           .COUT(co_mult_32u_32u_0_12_2), .S0(product_31__N_2324[9]), .S1(product_31__N_2324[10])) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(n41428), .B(store_m), .C(LM32D_CYC_O), 
         .D(n41512), .Z(w_clk_cpu_enable_623)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1676[29:48])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h0400;
    MULT2 mult_32u_32u_0_mult_0_3 (.A0(muliplicand[6]), .A1(muliplicand[7]), 
          .A2(muliplicand[7]), .A3(muliplicand[8]), .B0(operand_1_x[1]), 
          .B1(operand_1_x[0]), .B2(operand_1_x[1]), .B3(operand_1_x[0]), 
          .CI(mco_2), .CO(mco_3), .P0(mult_32u_32u_0_pp_0_7), .P1(mult_32u_32u_0_pp_0_8)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B Cadd_mult_32u_32u_0_12_1 (.A0(GND_net), .A1(s_mult_32u_32u_0_8_8), 
           .B0(GND_net), .B1(mult_32u_32u_0_pp_4_8), .CI(GND_net), .COUT(co_mult_32u_32u_0_12_1), 
           .S1(product_31__N_2324[8])) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_0_2 (.A0(muliplicand[4]), .A1(muliplicand[5]), 
          .A2(muliplicand[5]), .A3(muliplicand[6]), .B0(operand_1_x[1]), 
          .B1(operand_1_x[0]), .B2(operand_1_x[1]), .B3(operand_1_x[0]), 
          .CI(mco_1), .CO(mco_2), .P0(mult_32u_32u_0_pp_0_5), .P1(mult_32u_32u_0_pp_0_6)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    MULT2 mult_32u_32u_0_mult_0_1 (.A0(muliplicand[2]), .A1(muliplicand[3]), 
          .A2(muliplicand[3]), .A3(muliplicand[4]), .B0(operand_1_x[1]), 
          .B1(operand_1_x[0]), .B2(operand_1_x[1]), .B3(operand_1_x[0]), 
          .CI(mco), .CO(mco_1), .P0(mult_32u_32u_0_pp_0_3), .P1(mult_32u_32u_0_pp_0_4)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    LUT4 i1_2_lut_2_lut (.A(n41428), .B(store_m), .Z(n46)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1676[29:48])
    defparam i1_2_lut_2_lut.init = 16'h4444;
    MULT2 mult_32u_32u_0_mult_0_0 (.A0(muliplicand[0]), .A1(muliplicand[1]), 
          .A2(muliplicand[1]), .A3(muliplicand[2]), .B0(operand_1_x[1]), 
          .B1(operand_1_x[0]), .B2(operand_1_x[1]), .B3(operand_1_x[0]), 
          .CI(mult_32u_32u_0_cin_lr_0), .CO(mco), .P0(product_31__N_2324[1]), 
          .P1(mult_32u_32u_0_pp_0_2)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    LUT4 i20144_2_lut_2_lut (.A(n41428), .B(reset_exception), .Z(n22524)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1676[29:48])
    defparam i20144_2_lut_2_lut.init = 16'h4444;
    LUT4 i23498_3_lut_3_lut (.A(n41428), .B(\size_x[1] ), .C(\condition_x[0] ), 
         .Z(n26122)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1676[29:48])
    defparam i23498_3_lut_3_lut.init = 16'h1010;
    LUT4 i2_3_lut_4_lut_4_lut (.A(n41428), .B(n41513), .C(data_bus_error_exception), 
         .D(n41512), .Z(memop_pc_w_31__N_1219)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(1676[29:48])
    defparam i2_3_lut_4_lut_4_lut.init = 16'h0400;
    FADD2B t_mult_32u_32u_0_add_14_9 (.A0(s_mult_32u_32u_0_12_31), .A1(s_mult_32u_32u_0_12_32), 
           .B0(s_mult_32u_32u_0_13_31), .B1(s_mult_32u_32u_0_13_32), .CI(co_t_mult_32u_32u_0_14_8), 
           .S0(product_31__N_2324[31])) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B t_mult_32u_32u_0_add_14_8 (.A0(s_mult_32u_32u_0_12_29), .A1(s_mult_32u_32u_0_12_30), 
           .B0(s_mult_32u_32u_0_13_29), .B1(s_mult_32u_32u_0_13_30), .CI(co_t_mult_32u_32u_0_14_7), 
           .COUT(co_t_mult_32u_32u_0_14_8), .S0(product_31__N_2324[29]), 
           .S1(product_31__N_2324[30])) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B t_mult_32u_32u_0_add_14_7 (.A0(s_mult_32u_32u_0_12_27), .A1(s_mult_32u_32u_0_12_28), 
           .B0(s_mult_32u_32u_0_13_27), .B1(s_mult_32u_32u_0_13_28), .CI(co_t_mult_32u_32u_0_14_6), 
           .COUT(co_t_mult_32u_32u_0_14_7), .S0(product_31__N_2324[27]), 
           .S1(product_31__N_2324[28])) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B t_mult_32u_32u_0_add_14_6 (.A0(s_mult_32u_32u_0_12_25), .A1(s_mult_32u_32u_0_12_26), 
           .B0(s_mult_32u_32u_0_13_25), .B1(s_mult_32u_32u_0_13_26), .CI(co_t_mult_32u_32u_0_14_5), 
           .COUT(co_t_mult_32u_32u_0_14_6), .S0(product_31__N_2324[25]), 
           .S1(product_31__N_2324[26])) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B t_mult_32u_32u_0_add_14_5 (.A0(s_mult_32u_32u_0_12_23), .A1(s_mult_32u_32u_0_12_24), 
           .B0(s_mult_32u_32u_0_10_23), .B1(s_mult_32u_32u_0_13_24), .CI(co_t_mult_32u_32u_0_14_4), 
           .COUT(co_t_mult_32u_32u_0_14_5), .S0(product_31__N_2324[23]), 
           .S1(product_31__N_2324[24])) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B t_mult_32u_32u_0_add_14_4 (.A0(s_mult_32u_32u_0_12_21), .A1(s_mult_32u_32u_0_12_22), 
           .B0(s_mult_32u_32u_0_10_21), .B1(s_mult_32u_32u_0_10_22), .CI(co_t_mult_32u_32u_0_14_3), 
           .COUT(co_t_mult_32u_32u_0_14_4), .S0(product_31__N_2324[21]), 
           .S1(product_31__N_2324[22])) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B t_mult_32u_32u_0_add_14_3 (.A0(s_mult_32u_32u_0_12_19), .A1(s_mult_32u_32u_0_12_20), 
           .B0(s_mult_32u_32u_0_4_19), .B1(s_mult_32u_32u_0_10_20), .CI(co_t_mult_32u_32u_0_14_2), 
           .COUT(co_t_mult_32u_32u_0_14_3), .S0(product_31__N_2324[19]), 
           .S1(product_31__N_2324[20])) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B t_mult_32u_32u_0_add_14_2 (.A0(s_mult_32u_32u_0_12_17), .A1(s_mult_32u_32u_0_12_18), 
           .B0(mult_32u_32u_0_pp_8_17), .B1(s_mult_32u_32u_0_4_18), .CI(co_t_mult_32u_32u_0_14_1), 
           .COUT(co_t_mult_32u_32u_0_14_2), .S0(product_31__N_2324[17]), 
           .S1(product_31__N_2324[18])) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B Cadd_t_mult_32u_32u_0_14_1 (.A0(GND_net), .A1(s_mult_32u_32u_0_12_16), 
           .B0(GND_net), .B1(mult_32u_32u_0_pp_8_16), .CI(GND_net), .COUT(co_t_mult_32u_32u_0_14_1), 
           .S1(product_31__N_2324[16])) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_3_10 (.A0(mult_32u_32u_0_pp_6_31), .A1(mult_32u_32u_0_pp_6_32), 
           .B0(mult_32u_32u_0_pp_7_31), .B1(mult_32u_32u_0_pp_7_32), .CI(co_mult_32u_32u_0_3_9), 
           .S0(s_mult_32u_32u_0_3_31), .S1(s_mult_32u_32u_0_3_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_3_9 (.A0(mult_32u_32u_0_pp_6_29), .A1(mult_32u_32u_0_pp_6_30), 
           .B0(mult_32u_32u_0_pp_7_29), .B1(mult_32u_32u_0_pp_7_30), .CI(co_mult_32u_32u_0_3_8), 
           .COUT(co_mult_32u_32u_0_3_9), .S0(s_mult_32u_32u_0_3_29), .S1(s_mult_32u_32u_0_3_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_3_8 (.A0(mult_32u_32u_0_pp_6_27), .A1(mult_32u_32u_0_pp_6_28), 
           .B0(mult_32u_32u_0_pp_7_27), .B1(mult_32u_32u_0_pp_7_28), .CI(co_mult_32u_32u_0_3_7), 
           .COUT(co_mult_32u_32u_0_3_8), .S0(s_mult_32u_32u_0_3_27), .S1(s_mult_32u_32u_0_3_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_3_7 (.A0(mult_32u_32u_0_pp_6_25), .A1(mult_32u_32u_0_pp_6_26), 
           .B0(mult_32u_32u_0_pp_7_25), .B1(mult_32u_32u_0_pp_7_26), .CI(co_mult_32u_32u_0_3_6), 
           .COUT(co_mult_32u_32u_0_3_7), .S0(s_mult_32u_32u_0_3_25), .S1(s_mult_32u_32u_0_3_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_3_6 (.A0(mult_32u_32u_0_pp_6_23), .A1(mult_32u_32u_0_pp_6_24), 
           .B0(mult_32u_32u_0_pp_7_23), .B1(mult_32u_32u_0_pp_7_24), .CI(co_mult_32u_32u_0_3_5), 
           .COUT(co_mult_32u_32u_0_3_6), .S0(s_mult_32u_32u_0_3_23), .S1(s_mult_32u_32u_0_3_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_3_5 (.A0(mult_32u_32u_0_pp_6_21), .A1(mult_32u_32u_0_pp_6_22), 
           .B0(mult_32u_32u_0_pp_7_21), .B1(mult_32u_32u_0_pp_7_22), .CI(co_mult_32u_32u_0_3_4), 
           .COUT(co_mult_32u_32u_0_3_5), .S0(s_mult_32u_32u_0_3_21), .S1(s_mult_32u_32u_0_3_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_3_4 (.A0(mult_32u_32u_0_pp_6_19), .A1(mult_32u_32u_0_pp_6_20), 
           .B0(mult_32u_32u_0_pp_7_19), .B1(mult_32u_32u_0_pp_7_20), .CI(co_mult_32u_32u_0_3_3), 
           .COUT(co_mult_32u_32u_0_3_4), .S0(s_mult_32u_32u_0_3_19), .S1(s_mult_32u_32u_0_3_20)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_3_3 (.A0(mult_32u_32u_0_pp_6_17), .A1(mult_32u_32u_0_pp_6_18), 
           .B0(mult_32u_32u_0_pp_7_17), .B1(mult_32u_32u_0_pp_7_18), .CI(co_mult_32u_32u_0_3_2), 
           .COUT(co_mult_32u_32u_0_3_3), .S0(s_mult_32u_32u_0_3_17), .S1(s_mult_32u_32u_0_3_18)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_3_2 (.A0(mult_32u_32u_0_pp_6_15), .A1(mult_32u_32u_0_pp_6_16), 
           .B0(mult_32u_32u_0_pp_7_15), .B1(mult_32u_32u_0_pp_7_16), .CI(co_mult_32u_32u_0_3_1), 
           .COUT(co_mult_32u_32u_0_3_2), .S0(s_mult_32u_32u_0_3_15), .S1(s_mult_32u_32u_0_3_16)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B Cadd_mult_32u_32u_0_3_1 (.A0(GND_net), .A1(mult_32u_32u_0_pp_6_14), 
           .B0(GND_net), .B1(mult_32u_32u_0_pp_7_14), .CI(GND_net), .COUT(co_mult_32u_32u_0_3_1), 
           .S1(s_mult_32u_32u_0_3_14)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_11_3 (.A0(s_mult_32u_32u_0_6_31), .A1(s_mult_32u_32u_0_6_32), 
           .B0(s_mult_32u_32u_0_7_31), .B1(s_mult_32u_32u_0_7_32), .CI(co_mult_32u_32u_0_11_2), 
           .S0(s_mult_32u_32u_0_11_31), .S1(s_mult_32u_32u_0_11_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_11_2 (.A0(s_mult_32u_32u_0_6_29), .A1(s_mult_32u_32u_0_6_30), 
           .B0(mult_32u_32u_0_pp_14_29), .B1(s_mult_32u_32u_0_7_30), .CI(co_mult_32u_32u_0_11_1), 
           .COUT(co_mult_32u_32u_0_11_2), .S0(s_mult_32u_32u_0_11_29), .S1(s_mult_32u_32u_0_11_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_2_12 (.A0(mult_32u_32u_0_pp_4_31), .A1(mult_32u_32u_0_pp_4_32), 
           .B0(mult_32u_32u_0_pp_5_31), .B1(mult_32u_32u_0_pp_5_32), .CI(co_mult_32u_32u_0_2_11), 
           .S0(s_mult_32u_32u_0_2_31), .S1(s_mult_32u_32u_0_2_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B Cadd_mult_32u_32u_0_11_1 (.A0(GND_net), .A1(s_mult_32u_32u_0_6_28), 
           .B0(GND_net), .B1(mult_32u_32u_0_pp_14_28), .CI(GND_net), .COUT(co_mult_32u_32u_0_11_1), 
           .S1(s_mult_32u_32u_0_11_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_2_11 (.A0(mult_32u_32u_0_pp_4_29), .A1(mult_32u_32u_0_pp_4_30), 
           .B0(mult_32u_32u_0_pp_5_29), .B1(mult_32u_32u_0_pp_5_30), .CI(co_mult_32u_32u_0_2_10), 
           .COUT(co_mult_32u_32u_0_2_11), .S0(s_mult_32u_32u_0_2_29), .S1(s_mult_32u_32u_0_2_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_2_10 (.A0(mult_32u_32u_0_pp_4_27), .A1(mult_32u_32u_0_pp_4_28), 
           .B0(mult_32u_32u_0_pp_5_27), .B1(mult_32u_32u_0_pp_5_28), .CI(co_mult_32u_32u_0_2_9), 
           .COUT(co_mult_32u_32u_0_2_10), .S0(s_mult_32u_32u_0_2_27), .S1(s_mult_32u_32u_0_2_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_2_9 (.A0(mult_32u_32u_0_pp_4_25), .A1(mult_32u_32u_0_pp_4_26), 
           .B0(mult_32u_32u_0_pp_5_25), .B1(mult_32u_32u_0_pp_5_26), .CI(co_mult_32u_32u_0_2_8), 
           .COUT(co_mult_32u_32u_0_2_9), .S0(s_mult_32u_32u_0_2_25), .S1(s_mult_32u_32u_0_2_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_2_8 (.A0(mult_32u_32u_0_pp_4_23), .A1(mult_32u_32u_0_pp_4_24), 
           .B0(mult_32u_32u_0_pp_5_23), .B1(mult_32u_32u_0_pp_5_24), .CI(co_mult_32u_32u_0_2_7), 
           .COUT(co_mult_32u_32u_0_2_8), .S0(s_mult_32u_32u_0_2_23), .S1(s_mult_32u_32u_0_2_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_2_7 (.A0(mult_32u_32u_0_pp_4_21), .A1(mult_32u_32u_0_pp_4_22), 
           .B0(mult_32u_32u_0_pp_5_21), .B1(mult_32u_32u_0_pp_5_22), .CI(co_mult_32u_32u_0_2_6), 
           .COUT(co_mult_32u_32u_0_2_7), .S0(s_mult_32u_32u_0_2_21), .S1(s_mult_32u_32u_0_2_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_2_6 (.A0(mult_32u_32u_0_pp_4_19), .A1(mult_32u_32u_0_pp_4_20), 
           .B0(mult_32u_32u_0_pp_5_19), .B1(mult_32u_32u_0_pp_5_20), .CI(co_mult_32u_32u_0_2_5), 
           .COUT(co_mult_32u_32u_0_2_6), .S0(s_mult_32u_32u_0_2_19), .S1(s_mult_32u_32u_0_2_20)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_2_5 (.A0(mult_32u_32u_0_pp_4_17), .A1(mult_32u_32u_0_pp_4_18), 
           .B0(mult_32u_32u_0_pp_5_17), .B1(mult_32u_32u_0_pp_5_18), .CI(co_mult_32u_32u_0_2_4), 
           .COUT(co_mult_32u_32u_0_2_5), .S0(s_mult_32u_32u_0_2_17), .S1(s_mult_32u_32u_0_2_18)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_2_4 (.A0(mult_32u_32u_0_pp_4_15), .A1(mult_32u_32u_0_pp_4_16), 
           .B0(mult_32u_32u_0_pp_5_15), .B1(mult_32u_32u_0_pp_5_16), .CI(co_mult_32u_32u_0_2_3), 
           .COUT(co_mult_32u_32u_0_2_4), .S0(s_mult_32u_32u_0_2_15), .S1(s_mult_32u_32u_0_2_16)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_2_3 (.A0(mult_32u_32u_0_pp_4_13), .A1(mult_32u_32u_0_pp_4_14), 
           .B0(mult_32u_32u_0_pp_5_13), .B1(mult_32u_32u_0_pp_5_14), .CI(co_mult_32u_32u_0_2_2), 
           .COUT(co_mult_32u_32u_0_2_3), .S0(s_mult_32u_32u_0_2_13), .S1(s_mult_32u_32u_0_2_14)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_10_7 (.A0(s_mult_32u_32u_0_4_31), .A1(s_mult_32u_32u_0_4_32), 
           .B0(s_mult_32u_32u_0_5_31), .B1(s_mult_32u_32u_0_5_32), .CI(co_mult_32u_32u_0_10_6), 
           .S0(s_mult_32u_32u_0_10_31), .S1(s_mult_32u_32u_0_10_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_10_6 (.A0(s_mult_32u_32u_0_4_29), .A1(s_mult_32u_32u_0_4_30), 
           .B0(s_mult_32u_32u_0_5_29), .B1(s_mult_32u_32u_0_5_30), .CI(co_mult_32u_32u_0_10_5), 
           .COUT(co_mult_32u_32u_0_10_6), .S0(s_mult_32u_32u_0_10_29), .S1(s_mult_32u_32u_0_10_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_10_5 (.A0(s_mult_32u_32u_0_4_27), .A1(s_mult_32u_32u_0_4_28), 
           .B0(s_mult_32u_32u_0_5_27), .B1(s_mult_32u_32u_0_5_28), .CI(co_mult_32u_32u_0_10_4), 
           .COUT(co_mult_32u_32u_0_10_5), .S0(s_mult_32u_32u_0_10_27), .S1(s_mult_32u_32u_0_10_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1P3AX product_i0_i0 (.D(product_31__N_2324[0]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(product[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i0.GSR = "ENABLED";
    FD1S3AX result_i0 (.D(product[0]), .CK(w_clk_cpu), .Q(multiplier_result_w[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i0.GSR = "ENABLED";
    FADD2B mult_32u_32u_0_add_2_2 (.A0(mult_32u_32u_0_pp_4_11), .A1(mult_32u_32u_0_pp_4_12), 
           .B0(mult_32u_32u_0_pp_5_11), .B1(mult_32u_32u_0_pp_5_12), .CI(co_mult_32u_32u_0_2_1), 
           .COUT(co_mult_32u_32u_0_2_2), .S0(s_mult_32u_32u_0_2_11), .S1(s_mult_32u_32u_0_2_12)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B Cadd_mult_32u_32u_0_2_1 (.A0(GND_net), .A1(mult_32u_32u_0_pp_4_10), 
           .B0(GND_net), .B1(mult_32u_32u_0_pp_5_10), .CI(GND_net), .COUT(co_mult_32u_32u_0_2_1), 
           .S1(s_mult_32u_32u_0_2_10)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_10_4 (.A0(s_mult_32u_32u_0_4_25), .A1(s_mult_32u_32u_0_4_26), 
           .B0(s_mult_32u_32u_0_5_25), .B1(s_mult_32u_32u_0_5_26), .CI(co_mult_32u_32u_0_10_3), 
           .COUT(co_mult_32u_32u_0_10_4), .S0(s_mult_32u_32u_0_10_25), .S1(s_mult_32u_32u_0_10_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_10_3 (.A0(s_mult_32u_32u_0_4_23), .A1(s_mult_32u_32u_0_4_24), 
           .B0(s_mult_32u_32u_0_5_23), .B1(s_mult_32u_32u_0_5_24), .CI(co_mult_32u_32u_0_10_2), 
           .COUT(co_mult_32u_32u_0_10_3), .S0(s_mult_32u_32u_0_10_23), .S1(s_mult_32u_32u_0_10_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_10_2 (.A0(s_mult_32u_32u_0_4_21), .A1(s_mult_32u_32u_0_4_22), 
           .B0(mult_32u_32u_0_pp_10_21), .B1(s_mult_32u_32u_0_5_22), .CI(co_mult_32u_32u_0_10_1), 
           .COUT(co_mult_32u_32u_0_10_2), .S0(s_mult_32u_32u_0_10_21), .S1(s_mult_32u_32u_0_10_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B Cadd_mult_32u_32u_0_10_1 (.A0(GND_net), .A1(s_mult_32u_32u_0_4_20), 
           .B0(GND_net), .B1(mult_32u_32u_0_pp_10_20), .CI(GND_net), .COUT(co_mult_32u_32u_0_10_1), 
           .S1(s_mult_32u_32u_0_10_20)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_1_14 (.A0(mult_32u_32u_0_pp_2_31), .A1(mult_32u_32u_0_pp_2_32), 
           .B0(mult_32u_32u_0_pp_3_31), .B1(mult_32u_32u_0_pp_3_32), .CI(co_mult_32u_32u_0_1_13), 
           .S0(s_mult_32u_32u_0_1_31), .S1(s_mult_32u_32u_0_1_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_1_13 (.A0(mult_32u_32u_0_pp_2_29), .A1(mult_32u_32u_0_pp_2_30), 
           .B0(mult_32u_32u_0_pp_3_29), .B1(mult_32u_32u_0_pp_3_30), .CI(co_mult_32u_32u_0_1_12), 
           .COUT(co_mult_32u_32u_0_1_13), .S0(s_mult_32u_32u_0_1_29), .S1(s_mult_32u_32u_0_1_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_1_12 (.A0(mult_32u_32u_0_pp_2_27), .A1(mult_32u_32u_0_pp_2_28), 
           .B0(mult_32u_32u_0_pp_3_27), .B1(mult_32u_32u_0_pp_3_28), .CI(co_mult_32u_32u_0_1_11), 
           .COUT(co_mult_32u_32u_0_1_12), .S0(s_mult_32u_32u_0_1_27), .S1(s_mult_32u_32u_0_1_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_1_11 (.A0(mult_32u_32u_0_pp_2_25), .A1(mult_32u_32u_0_pp_2_26), 
           .B0(mult_32u_32u_0_pp_3_25), .B1(mult_32u_32u_0_pp_3_26), .CI(co_mult_32u_32u_0_1_10), 
           .COUT(co_mult_32u_32u_0_1_11), .S0(s_mult_32u_32u_0_1_25), .S1(s_mult_32u_32u_0_1_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_1_10 (.A0(mult_32u_32u_0_pp_2_23), .A1(mult_32u_32u_0_pp_2_24), 
           .B0(mult_32u_32u_0_pp_3_23), .B1(mult_32u_32u_0_pp_3_24), .CI(co_mult_32u_32u_0_1_9), 
           .COUT(co_mult_32u_32u_0_1_10), .S0(s_mult_32u_32u_0_1_23), .S1(s_mult_32u_32u_0_1_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_1_9 (.A0(mult_32u_32u_0_pp_2_21), .A1(mult_32u_32u_0_pp_2_22), 
           .B0(mult_32u_32u_0_pp_3_21), .B1(mult_32u_32u_0_pp_3_22), .CI(co_mult_32u_32u_0_1_8), 
           .COUT(co_mult_32u_32u_0_1_9), .S0(s_mult_32u_32u_0_1_21), .S1(s_mult_32u_32u_0_1_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_1_8 (.A0(mult_32u_32u_0_pp_2_19), .A1(mult_32u_32u_0_pp_2_20), 
           .B0(mult_32u_32u_0_pp_3_19), .B1(mult_32u_32u_0_pp_3_20), .CI(co_mult_32u_32u_0_1_7), 
           .COUT(co_mult_32u_32u_0_1_8), .S0(s_mult_32u_32u_0_1_19), .S1(s_mult_32u_32u_0_1_20)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_9_11 (.A0(s_mult_32u_32u_0_2_31), .A1(s_mult_32u_32u_0_2_32), 
           .B0(s_mult_32u_32u_0_3_31), .B1(s_mult_32u_32u_0_3_32), .CI(co_mult_32u_32u_0_9_10), 
           .S0(s_mult_32u_32u_0_9_31), .S1(s_mult_32u_32u_0_9_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_9_10 (.A0(s_mult_32u_32u_0_2_29), .A1(s_mult_32u_32u_0_2_30), 
           .B0(s_mult_32u_32u_0_3_29), .B1(s_mult_32u_32u_0_3_30), .CI(co_mult_32u_32u_0_9_9), 
           .COUT(co_mult_32u_32u_0_9_10), .S0(s_mult_32u_32u_0_9_29), .S1(s_mult_32u_32u_0_9_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_1_7 (.A0(mult_32u_32u_0_pp_2_17), .A1(mult_32u_32u_0_pp_2_18), 
           .B0(mult_32u_32u_0_pp_3_17), .B1(mult_32u_32u_0_pp_3_18), .CI(co_mult_32u_32u_0_1_6), 
           .COUT(co_mult_32u_32u_0_1_7), .S0(s_mult_32u_32u_0_1_17), .S1(s_mult_32u_32u_0_1_18)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_1_6 (.A0(mult_32u_32u_0_pp_2_15), .A1(mult_32u_32u_0_pp_2_16), 
           .B0(mult_32u_32u_0_pp_3_15), .B1(mult_32u_32u_0_pp_3_16), .CI(co_mult_32u_32u_0_1_5), 
           .COUT(co_mult_32u_32u_0_1_6), .S0(s_mult_32u_32u_0_1_15), .S1(s_mult_32u_32u_0_1_16)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_1_5 (.A0(mult_32u_32u_0_pp_2_13), .A1(mult_32u_32u_0_pp_2_14), 
           .B0(mult_32u_32u_0_pp_3_13), .B1(mult_32u_32u_0_pp_3_14), .CI(co_mult_32u_32u_0_1_4), 
           .COUT(co_mult_32u_32u_0_1_5), .S0(s_mult_32u_32u_0_1_13), .S1(s_mult_32u_32u_0_1_14)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_1_4 (.A0(mult_32u_32u_0_pp_2_11), .A1(mult_32u_32u_0_pp_2_12), 
           .B0(mult_32u_32u_0_pp_3_11), .B1(mult_32u_32u_0_pp_3_12), .CI(co_mult_32u_32u_0_1_3), 
           .COUT(co_mult_32u_32u_0_1_4), .S0(s_mult_32u_32u_0_1_11), .S1(s_mult_32u_32u_0_1_12)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_1_3 (.A0(mult_32u_32u_0_pp_2_9), .A1(mult_32u_32u_0_pp_2_10), 
           .B0(mult_32u_32u_0_pp_3_9), .B1(mult_32u_32u_0_pp_3_10), .CI(co_mult_32u_32u_0_1_2), 
           .COUT(co_mult_32u_32u_0_1_3), .S0(s_mult_32u_32u_0_1_9), .S1(s_mult_32u_32u_0_1_10)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_1_2 (.A0(mult_32u_32u_0_pp_2_7), .A1(mult_32u_32u_0_pp_2_8), 
           .B0(mult_32u_32u_0_pp_3_7), .B1(mult_32u_32u_0_pp_3_8), .CI(co_mult_32u_32u_0_1_1), 
           .COUT(co_mult_32u_32u_0_1_2), .S0(s_mult_32u_32u_0_1_7), .S1(s_mult_32u_32u_0_1_8)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B Cadd_mult_32u_32u_0_1_1 (.A0(GND_net), .A1(mult_32u_32u_0_pp_2_6), 
           .B0(GND_net), .B1(mult_32u_32u_0_pp_3_6), .CI(GND_net), .COUT(co_mult_32u_32u_0_1_1), 
           .S1(s_mult_32u_32u_0_1_6)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_9_9 (.A0(s_mult_32u_32u_0_2_27), .A1(s_mult_32u_32u_0_2_28), 
           .B0(s_mult_32u_32u_0_3_27), .B1(s_mult_32u_32u_0_3_28), .CI(co_mult_32u_32u_0_9_8), 
           .COUT(co_mult_32u_32u_0_9_9), .S0(s_mult_32u_32u_0_9_27), .S1(s_mult_32u_32u_0_9_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_9_8 (.A0(s_mult_32u_32u_0_2_25), .A1(s_mult_32u_32u_0_2_26), 
           .B0(s_mult_32u_32u_0_3_25), .B1(s_mult_32u_32u_0_3_26), .CI(co_mult_32u_32u_0_9_7), 
           .COUT(co_mult_32u_32u_0_9_8), .S0(s_mult_32u_32u_0_9_25), .S1(s_mult_32u_32u_0_9_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_0_16 (.A0(mult_32u_32u_0_pp_0_31), .A1(mult_32u_32u_0_pp_0_32), 
           .B0(mult_32u_32u_0_pp_1_31), .B1(mult_32u_32u_0_pp_1_32), .CI(co_mult_32u_32u_0_0_15), 
           .S0(s_mult_32u_32u_0_0_31), .S1(s_mult_32u_32u_0_0_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_0_15 (.A0(mult_32u_32u_0_pp_0_29), .A1(mult_32u_32u_0_pp_0_30), 
           .B0(mult_32u_32u_0_pp_1_29), .B1(mult_32u_32u_0_pp_1_30), .CI(co_mult_32u_32u_0_0_14), 
           .COUT(co_mult_32u_32u_0_0_15), .S0(s_mult_32u_32u_0_0_29), .S1(s_mult_32u_32u_0_0_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_0_14 (.A0(mult_32u_32u_0_pp_0_27), .A1(mult_32u_32u_0_pp_0_28), 
           .B0(mult_32u_32u_0_pp_1_27), .B1(mult_32u_32u_0_pp_1_28), .CI(co_mult_32u_32u_0_0_13), 
           .COUT(co_mult_32u_32u_0_0_14), .S0(s_mult_32u_32u_0_0_27), .S1(s_mult_32u_32u_0_0_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_0_13 (.A0(mult_32u_32u_0_pp_0_25), .A1(mult_32u_32u_0_pp_0_26), 
           .B0(mult_32u_32u_0_pp_1_25), .B1(mult_32u_32u_0_pp_1_26), .CI(co_mult_32u_32u_0_0_12), 
           .COUT(co_mult_32u_32u_0_0_13), .S0(s_mult_32u_32u_0_0_25), .S1(s_mult_32u_32u_0_0_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_0_12 (.A0(mult_32u_32u_0_pp_0_23), .A1(mult_32u_32u_0_pp_0_24), 
           .B0(mult_32u_32u_0_pp_1_23), .B1(mult_32u_32u_0_pp_1_24), .CI(co_mult_32u_32u_0_0_11), 
           .COUT(co_mult_32u_32u_0_0_12), .S0(s_mult_32u_32u_0_0_23), .S1(s_mult_32u_32u_0_0_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_0_11 (.A0(mult_32u_32u_0_pp_0_21), .A1(mult_32u_32u_0_pp_0_22), 
           .B0(mult_32u_32u_0_pp_1_21), .B1(mult_32u_32u_0_pp_1_22), .CI(co_mult_32u_32u_0_0_10), 
           .COUT(co_mult_32u_32u_0_0_11), .S0(s_mult_32u_32u_0_0_21), .S1(s_mult_32u_32u_0_0_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_9_7 (.A0(s_mult_32u_32u_0_2_23), .A1(s_mult_32u_32u_0_2_24), 
           .B0(s_mult_32u_32u_0_3_23), .B1(s_mult_32u_32u_0_3_24), .CI(co_mult_32u_32u_0_9_6), 
           .COUT(co_mult_32u_32u_0_9_7), .S0(s_mult_32u_32u_0_9_23), .S1(s_mult_32u_32u_0_9_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_0_10 (.A0(mult_32u_32u_0_pp_0_19), .A1(mult_32u_32u_0_pp_0_20), 
           .B0(mult_32u_32u_0_pp_1_19), .B1(mult_32u_32u_0_pp_1_20), .CI(co_mult_32u_32u_0_0_9), 
           .COUT(co_mult_32u_32u_0_0_10), .S0(s_mult_32u_32u_0_0_19), .S1(s_mult_32u_32u_0_0_20)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_0_9 (.A0(mult_32u_32u_0_pp_0_17), .A1(mult_32u_32u_0_pp_0_18), 
           .B0(mult_32u_32u_0_pp_1_17), .B1(mult_32u_32u_0_pp_1_18), .CI(co_mult_32u_32u_0_0_8), 
           .COUT(co_mult_32u_32u_0_0_9), .S0(s_mult_32u_32u_0_0_17), .S1(s_mult_32u_32u_0_0_18)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_9_6 (.A0(s_mult_32u_32u_0_2_21), .A1(s_mult_32u_32u_0_2_22), 
           .B0(s_mult_32u_32u_0_3_21), .B1(s_mult_32u_32u_0_3_22), .CI(co_mult_32u_32u_0_9_5), 
           .COUT(co_mult_32u_32u_0_9_6), .S0(s_mult_32u_32u_0_9_21), .S1(s_mult_32u_32u_0_9_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_0_8 (.A0(mult_32u_32u_0_pp_0_15), .A1(mult_32u_32u_0_pp_0_16), 
           .B0(mult_32u_32u_0_pp_1_15), .B1(mult_32u_32u_0_pp_1_16), .CI(co_mult_32u_32u_0_0_7), 
           .COUT(co_mult_32u_32u_0_0_8), .S0(s_mult_32u_32u_0_0_15), .S1(s_mult_32u_32u_0_0_16)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_9_5 (.A0(s_mult_32u_32u_0_2_19), .A1(s_mult_32u_32u_0_2_20), 
           .B0(s_mult_32u_32u_0_3_19), .B1(s_mult_32u_32u_0_3_20), .CI(co_mult_32u_32u_0_9_4), 
           .COUT(co_mult_32u_32u_0_9_5), .S0(s_mult_32u_32u_0_9_19), .S1(s_mult_32u_32u_0_9_20)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    AND2 AND2_t11 (.A(muliplicand[0]), .B(operand_1_x[8]), .Z(mult_32u_32u_0_pp_4_8)) /* synthesis syn_instantiated=1 */ ;   // mult_32u_32u.v(1662[10:66])
    FADD2B mult_32u_32u_0_add_0_7 (.A0(mult_32u_32u_0_pp_0_13), .A1(mult_32u_32u_0_pp_0_14), 
           .B0(mult_32u_32u_0_pp_1_13), .B1(mult_32u_32u_0_pp_1_14), .CI(co_mult_32u_32u_0_0_6), 
           .COUT(co_mult_32u_32u_0_0_7), .S0(s_mult_32u_32u_0_0_13), .S1(s_mult_32u_32u_0_0_14)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_0_6 (.A0(mult_32u_32u_0_pp_0_11), .A1(mult_32u_32u_0_pp_0_12), 
           .B0(mult_32u_32u_0_pp_1_11), .B1(mult_32u_32u_0_pp_1_12), .CI(co_mult_32u_32u_0_0_5), 
           .COUT(co_mult_32u_32u_0_0_6), .S0(s_mult_32u_32u_0_0_11), .S1(s_mult_32u_32u_0_0_12)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_0_5 (.A0(mult_32u_32u_0_pp_0_9), .A1(mult_32u_32u_0_pp_0_10), 
           .B0(mult_32u_32u_0_pp_1_9), .B1(mult_32u_32u_0_pp_1_10), .CI(co_mult_32u_32u_0_0_4), 
           .COUT(co_mult_32u_32u_0_0_5), .S0(s_mult_32u_32u_0_0_9), .S1(s_mult_32u_32u_0_0_10)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_0_4 (.A0(mult_32u_32u_0_pp_0_7), .A1(mult_32u_32u_0_pp_0_8), 
           .B0(mult_32u_32u_0_pp_1_7), .B1(mult_32u_32u_0_pp_1_8), .CI(co_mult_32u_32u_0_0_3), 
           .COUT(co_mult_32u_32u_0_0_4), .S0(s_mult_32u_32u_0_0_7), .S1(s_mult_32u_32u_0_0_8)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1S3AX result_i14 (.D(product[14]), .CK(w_clk_cpu), .Q(multiplier_result_w[14])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i14.GSR = "ENABLED";
    FADD2B mult_32u_32u_0_add_0_3 (.A0(mult_32u_32u_0_pp_0_5), .A1(mult_32u_32u_0_pp_0_6), 
           .B0(mult_32u_32u_0_pp_1_5), .B1(mult_32u_32u_0_pp_1_6), .CI(co_mult_32u_32u_0_0_2), 
           .COUT(co_mult_32u_32u_0_0_3), .S0(s_mult_32u_32u_0_0_5), .S1(s_mult_32u_32u_0_0_6)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_0_2 (.A0(mult_32u_32u_0_pp_0_3), .A1(mult_32u_32u_0_pp_0_4), 
           .B0(mult_32u_32u_0_pp_1_3), .B1(mult_32u_32u_0_pp_1_4), .CI(co_mult_32u_32u_0_0_1), 
           .COUT(co_mult_32u_32u_0_0_2), .S0(product_31__N_2324[3]), .S1(s_mult_32u_32u_0_0_4)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B Cadd_mult_32u_32u_0_0_1 (.A0(GND_net), .A1(mult_32u_32u_0_pp_0_2), 
           .B0(GND_net), .B1(mult_32u_32u_0_pp_1_2), .CI(GND_net), .COUT(co_mult_32u_32u_0_0_1), 
           .S1(product_31__N_2324[2])) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1S3AX result_i13 (.D(product[13]), .CK(w_clk_cpu), .Q(multiplier_result_w[13])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i13.GSR = "ENABLED";
    FADD2B mult_32u_32u_0_cin_lr_add_30 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_32u_32u_0_cin_lr_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_cin_lr_add_28 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_32u_32u_0_cin_lr_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_9_4 (.A0(s_mult_32u_32u_0_2_17), .A1(s_mult_32u_32u_0_2_18), 
           .B0(s_mult_32u_32u_0_3_17), .B1(s_mult_32u_32u_0_3_18), .CI(co_mult_32u_32u_0_9_3), 
           .COUT(co_mult_32u_32u_0_9_4), .S0(s_mult_32u_32u_0_9_17), .S1(s_mult_32u_32u_0_9_18)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_9_3 (.A0(s_mult_32u_32u_0_2_15), .A1(s_mult_32u_32u_0_2_16), 
           .B0(s_mult_32u_32u_0_3_15), .B1(s_mult_32u_32u_0_3_16), .CI(co_mult_32u_32u_0_9_2), 
           .COUT(co_mult_32u_32u_0_9_3), .S0(s_mult_32u_32u_0_9_15), .S1(s_mult_32u_32u_0_9_16)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1S3AX result_i12 (.D(product[12]), .CK(w_clk_cpu), .Q(multiplier_result_w[12])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i12.GSR = "ENABLED";
    FADD2B mult_32u_32u_0_cin_lr_add_26 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_32u_32u_0_cin_lr_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_cin_lr_add_24 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_32u_32u_0_cin_lr_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_9_2 (.A0(s_mult_32u_32u_0_2_13), .A1(s_mult_32u_32u_0_2_14), 
           .B0(mult_32u_32u_0_pp_6_13), .B1(s_mult_32u_32u_0_3_14), .CI(co_mult_32u_32u_0_9_1), 
           .COUT(co_mult_32u_32u_0_9_2), .S0(s_mult_32u_32u_0_9_13), .S1(s_mult_32u_32u_0_9_14)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1S3AX result_i11 (.D(product[11]), .CK(w_clk_cpu), .Q(multiplier_result_w[11])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i11.GSR = "ENABLED";
    FADD2B mult_32u_32u_0_cin_lr_add_22 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_32u_32u_0_cin_lr_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_cin_lr_add_20 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_32u_32u_0_cin_lr_20)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1S3AX result_i10 (.D(product[10]), .CK(w_clk_cpu), .Q(multiplier_result_w[10])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i10.GSR = "ENABLED";
    FADD2B mult_32u_32u_0_cin_lr_add_18 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_32u_32u_0_cin_lr_18)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_cin_lr_add_16 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_32u_32u_0_cin_lr_16)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_cin_lr_add_14 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_32u_32u_0_cin_lr_14)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_cin_lr_add_12 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_32u_32u_0_cin_lr_12)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_cin_lr_add_10 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_32u_32u_0_cin_lr_10)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1S3AX result_i9 (.D(product[9]), .CK(w_clk_cpu), .Q(multiplier_result_w[9])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i9.GSR = "ENABLED";
    FADD2B Cadd_mult_32u_32u_0_9_1 (.A0(GND_net), .A1(s_mult_32u_32u_0_2_12), 
           .B0(GND_net), .B1(mult_32u_32u_0_pp_6_12), .CI(GND_net), .COUT(co_mult_32u_32u_0_9_1), 
           .S1(s_mult_32u_32u_0_9_12)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_cin_lr_add_8 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_32u_32u_0_cin_lr_8)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1S3AX result_i8 (.D(product[8]), .CK(w_clk_cpu), .Q(multiplier_result_w[8])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i8.GSR = "ENABLED";
    FADD2B mult_32u_32u_0_cin_lr_add_6 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_32u_32u_0_cin_lr_6)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_cin_lr_add_4 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_32u_32u_0_cin_lr_4)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_cin_lr_add_2 (.A0(GND_net), .A1(GND_net), .B0(GND_net), 
           .B1(GND_net), .CI(GND_net), .COUT(mult_32u_32u_0_cin_lr_2)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    AND2 AND2_t15 (.A(muliplicand[0]), .B(operand_1_x[0]), .Z(product_31__N_2324[0])) /* synthesis syn_instantiated=1 */ ;   // mult_32u_32u.v(1654[10:66])
    AND2 AND2_t14 (.A(muliplicand[0]), .B(operand_1_x[2]), .Z(mult_32u_32u_0_pp_1_2)) /* synthesis syn_instantiated=1 */ ;   // mult_32u_32u.v(1656[10:66])
    AND2 AND2_t13 (.A(muliplicand[0]), .B(operand_1_x[4]), .Z(mult_32u_32u_0_pp_2_4)) /* synthesis syn_instantiated=1 */ ;   // mult_32u_32u.v(1658[10:66])
    AND2 AND2_t12 (.A(muliplicand[0]), .B(operand_1_x[6]), .Z(mult_32u_32u_0_pp_3_6)) /* synthesis syn_instantiated=1 */ ;   // mult_32u_32u.v(1660[10:66])
    FD1S3AX result_i7 (.D(product[7]), .CK(w_clk_cpu), .Q(multiplier_result_w[7])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i7.GSR = "ENABLED";
    FD1S3AX result_i6 (.D(product[6]), .CK(w_clk_cpu), .Q(multiplier_result_w[6])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i6.GSR = "ENABLED";
    FD1S3AX result_i5 (.D(product[5]), .CK(w_clk_cpu), .Q(multiplier_result_w[5])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i5.GSR = "ENABLED";
    FD1S3AX result_i4 (.D(product[4]), .CK(w_clk_cpu), .Q(multiplier_result_w[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i4.GSR = "ENABLED";
    FADD2B mult_32u_32u_0_add_8_15 (.A0(s_mult_32u_32u_0_0_31), .A1(s_mult_32u_32u_0_0_32), 
           .B0(s_mult_32u_32u_0_1_31), .B1(s_mult_32u_32u_0_1_32), .CI(co_mult_32u_32u_0_8_14), 
           .S0(s_mult_32u_32u_0_8_31), .S1(s_mult_32u_32u_0_8_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_8_14 (.A0(s_mult_32u_32u_0_0_29), .A1(s_mult_32u_32u_0_0_30), 
           .B0(s_mult_32u_32u_0_1_29), .B1(s_mult_32u_32u_0_1_30), .CI(co_mult_32u_32u_0_8_13), 
           .COUT(co_mult_32u_32u_0_8_14), .S0(s_mult_32u_32u_0_8_29), .S1(s_mult_32u_32u_0_8_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1S3AX result_i3 (.D(product[3]), .CK(w_clk_cpu), .Q(multiplier_result_w[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i3.GSR = "ENABLED";
    FD1S3AX result_i2 (.D(product[2]), .CK(w_clk_cpu), .Q(multiplier_result_w[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i2.GSR = "ENABLED";
    FD1S3AX result_i1 (.D(product[1]), .CK(w_clk_cpu), .Q(multiplier_result_w[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i1.GSR = "ENABLED";
    FADD2B mult_32u_32u_0_add_8_13 (.A0(s_mult_32u_32u_0_0_27), .A1(s_mult_32u_32u_0_0_28), 
           .B0(s_mult_32u_32u_0_1_27), .B1(s_mult_32u_32u_0_1_28), .CI(co_mult_32u_32u_0_8_12), 
           .COUT(co_mult_32u_32u_0_8_13), .S0(s_mult_32u_32u_0_8_27), .S1(s_mult_32u_32u_0_8_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_8_12 (.A0(s_mult_32u_32u_0_0_25), .A1(s_mult_32u_32u_0_0_26), 
           .B0(s_mult_32u_32u_0_1_25), .B1(s_mult_32u_32u_0_1_26), .CI(co_mult_32u_32u_0_8_11), 
           .COUT(co_mult_32u_32u_0_8_12), .S0(s_mult_32u_32u_0_8_25), .S1(s_mult_32u_32u_0_8_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_8_11 (.A0(s_mult_32u_32u_0_0_23), .A1(s_mult_32u_32u_0_0_24), 
           .B0(s_mult_32u_32u_0_1_23), .B1(s_mult_32u_32u_0_1_24), .CI(co_mult_32u_32u_0_8_10), 
           .COUT(co_mult_32u_32u_0_8_11), .S0(s_mult_32u_32u_0_8_23), .S1(s_mult_32u_32u_0_8_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_8_10 (.A0(s_mult_32u_32u_0_0_21), .A1(s_mult_32u_32u_0_0_22), 
           .B0(s_mult_32u_32u_0_1_21), .B1(s_mult_32u_32u_0_1_22), .CI(co_mult_32u_32u_0_8_9), 
           .COUT(co_mult_32u_32u_0_8_10), .S0(s_mult_32u_32u_0_8_21), .S1(s_mult_32u_32u_0_8_22)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_8_9 (.A0(s_mult_32u_32u_0_0_19), .A1(s_mult_32u_32u_0_0_20), 
           .B0(s_mult_32u_32u_0_1_19), .B1(s_mult_32u_32u_0_1_20), .CI(co_mult_32u_32u_0_8_8), 
           .COUT(co_mult_32u_32u_0_8_9), .S0(s_mult_32u_32u_0_8_19), .S1(s_mult_32u_32u_0_8_20)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_8_8 (.A0(s_mult_32u_32u_0_0_17), .A1(s_mult_32u_32u_0_0_18), 
           .B0(s_mult_32u_32u_0_1_17), .B1(s_mult_32u_32u_0_1_18), .CI(co_mult_32u_32u_0_8_7), 
           .COUT(co_mult_32u_32u_0_8_8), .S0(s_mult_32u_32u_0_8_17), .S1(s_mult_32u_32u_0_8_18)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_8_7 (.A0(s_mult_32u_32u_0_0_15), .A1(s_mult_32u_32u_0_0_16), 
           .B0(s_mult_32u_32u_0_1_15), .B1(s_mult_32u_32u_0_1_16), .CI(co_mult_32u_32u_0_8_6), 
           .COUT(co_mult_32u_32u_0_8_7), .S0(s_mult_32u_32u_0_8_15), .S1(s_mult_32u_32u_0_8_16)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_8_6 (.A0(s_mult_32u_32u_0_0_13), .A1(s_mult_32u_32u_0_0_14), 
           .B0(s_mult_32u_32u_0_1_13), .B1(s_mult_32u_32u_0_1_14), .CI(co_mult_32u_32u_0_8_5), 
           .COUT(co_mult_32u_32u_0_8_6), .S0(s_mult_32u_32u_0_8_13), .S1(s_mult_32u_32u_0_8_14)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_8_5 (.A0(s_mult_32u_32u_0_0_11), .A1(s_mult_32u_32u_0_0_12), 
           .B0(s_mult_32u_32u_0_1_11), .B1(s_mult_32u_32u_0_1_12), .CI(co_mult_32u_32u_0_8_4), 
           .COUT(co_mult_32u_32u_0_8_5), .S0(s_mult_32u_32u_0_8_11), .S1(s_mult_32u_32u_0_8_12)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_8_4 (.A0(s_mult_32u_32u_0_0_9), .A1(s_mult_32u_32u_0_0_10), 
           .B0(s_mult_32u_32u_0_1_9), .B1(s_mult_32u_32u_0_1_10), .CI(co_mult_32u_32u_0_8_3), 
           .COUT(co_mult_32u_32u_0_8_4), .S0(s_mult_32u_32u_0_8_9), .S1(s_mult_32u_32u_0_8_10)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_8_3 (.A0(s_mult_32u_32u_0_0_7), .A1(s_mult_32u_32u_0_0_8), 
           .B0(s_mult_32u_32u_0_1_7), .B1(s_mult_32u_32u_0_1_8), .CI(co_mult_32u_32u_0_8_2), 
           .COUT(co_mult_32u_32u_0_8_3), .S0(product_31__N_2324[7]), .S1(s_mult_32u_32u_0_8_8)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_8_2 (.A0(s_mult_32u_32u_0_0_5), .A1(s_mult_32u_32u_0_0_6), 
           .B0(mult_32u_32u_0_pp_2_5), .B1(s_mult_32u_32u_0_1_6), .CI(co_mult_32u_32u_0_8_1), 
           .COUT(co_mult_32u_32u_0_8_2), .S0(product_31__N_2324[5]), .S1(product_31__N_2324[6])) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B Cadd_mult_32u_32u_0_8_1 (.A0(GND_net), .A1(s_mult_32u_32u_0_0_4), 
           .B0(GND_net), .B1(mult_32u_32u_0_pp_2_4), .CI(GND_net), .COUT(co_mult_32u_32u_0_8_1), 
           .S1(product_31__N_2324[4])) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1P3AX product_i0_i31 (.D(product_31__N_2324[31]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(product[31])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i31.GSR = "ENABLED";
    FD1P3AX product_i0_i30 (.D(product_31__N_2324[30]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(product[30])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i30.GSR = "ENABLED";
    FD1P3AX product_i0_i29 (.D(product_31__N_2324[29]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(product[29])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i29.GSR = "ENABLED";
    FD1P3AX product_i0_i28 (.D(product_31__N_2324[28]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(product[28])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i28.GSR = "ENABLED";
    FD1P3AX product_i0_i27 (.D(product_31__N_2324[27]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(product[27])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i27.GSR = "ENABLED";
    FD1P3AX product_i0_i26 (.D(product_31__N_2324[26]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(product[26])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i26.GSR = "ENABLED";
    FD1P3IX muliplicand_i0_i1 (.D(\bypass_data_0[1] ), .SP(w_clk_cpu_enable_984), 
            .CD(n26142), .CK(w_clk_cpu), .Q(muliplicand[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i1.GSR = "ENABLED";
    FD1P3AX product_i0_i25 (.D(product_31__N_2324[25]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(product[25])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i25.GSR = "ENABLED";
    FD1P3AX product_i0_i24 (.D(product_31__N_2324[24]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(product[24])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i24.GSR = "ENABLED";
    FD1P3AX product_i0_i23 (.D(product_31__N_2324[23]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(product[23])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i23.GSR = "ENABLED";
    FD1P3AX product_i0_i22 (.D(product_31__N_2324[22]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(product[22])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i22.GSR = "ENABLED";
    FD1P3AX product_i0_i21 (.D(product_31__N_2324[21]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(product[21])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i21.GSR = "ENABLED";
    FD1P3AX product_i0_i20 (.D(product_31__N_2324[20]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(product[20])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i20.GSR = "ENABLED";
    FD1P3AX product_i0_i19 (.D(product_31__N_2324[19]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(product[19])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i19.GSR = "ENABLED";
    FD1P3AX product_i0_i18 (.D(product_31__N_2324[18]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(product[18])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i18.GSR = "ENABLED";
    FD1P3IX muliplicand_i0_i0 (.D(\bypass_data_0[0] ), .SP(w_clk_cpu_enable_984), 
            .CD(n26142), .CK(w_clk_cpu), .Q(muliplicand[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i0.GSR = "ENABLED";
    FD1P3AX product_i0_i17 (.D(product_31__N_2324[17]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(product[17])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i17.GSR = "ENABLED";
    FD1P3AX product_i0_i16 (.D(product_31__N_2324[16]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(product[16])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i16.GSR = "ENABLED";
    FD1P3AX product_i0_i15 (.D(product_31__N_2324[15]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(product[15])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i15.GSR = "ENABLED";
    FD1P3AX product_i0_i14 (.D(product_31__N_2324[14]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(product[14])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i14.GSR = "ENABLED";
    FD1P3AX product_i0_i13 (.D(product_31__N_2324[13]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(product[13])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i13.GSR = "ENABLED";
    FD1P3AX product_i0_i12 (.D(product_31__N_2324[12]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(product[12])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i12.GSR = "ENABLED";
    FD1P3AX product_i0_i11 (.D(product_31__N_2324[11]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(product[11])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i11.GSR = "ENABLED";
    FD1P3AX product_i0_i10 (.D(product_31__N_2324[10]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(product[10])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i10.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i31 (.D(\d_result_0[31] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[31])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i31.GSR = "ENABLED";
    FD1P3AX product_i0_i9 (.D(product_31__N_2324[9]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(product[9])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i9.GSR = "ENABLED";
    FD1P3AX product_i0_i8 (.D(product_31__N_2324[8]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(product[8])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i8.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i30 (.D(\d_result_0[30] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[30])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i30.GSR = "ENABLED";
    FADD2B mult_32u_32u_0_add_7_2 (.A0(mult_32u_32u_0_pp_14_31), .A1(mult_32u_32u_0_pp_14_32), 
           .B0(mult_32u_32u_0_pp_15_31), .B1(mult_32u_32u_0_pp_15_32), .CI(co_mult_32u_32u_0_7_1), 
           .S0(s_mult_32u_32u_0_7_31), .S1(s_mult_32u_32u_0_7_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1P3AX product_i0_i7 (.D(product_31__N_2324[7]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(product[7])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i7.GSR = "ENABLED";
    FD1P3AX product_i0_i6 (.D(product_31__N_2324[6]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(product[6])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i6.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i29 (.D(\d_result_0[29] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[29])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i29.GSR = "ENABLED";
    FADD2B Cadd_mult_32u_32u_0_7_1 (.A0(GND_net), .A1(mult_32u_32u_0_pp_14_30), 
           .B0(GND_net), .B1(mult_32u_32u_0_pp_15_30), .CI(GND_net), .COUT(co_mult_32u_32u_0_7_1), 
           .S1(s_mult_32u_32u_0_7_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1P3AX product_i0_i5 (.D(product_31__N_2324[5]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(product[5])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i5.GSR = "ENABLED";
    FD1P3AX product_i0_i4 (.D(product_31__N_2324[4]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(product[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i4.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i28 (.D(\d_result_0[28] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[28])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i28.GSR = "ENABLED";
    FD1P3AX product_i0_i3 (.D(product_31__N_2324[3]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(product[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i3.GSR = "ENABLED";
    FD1P3AX product_i0_i2 (.D(product_31__N_2324[2]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(product[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i2.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i27 (.D(\d_result_0[27] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[27])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i27.GSR = "ENABLED";
    FD1P3AX product_i0_i1 (.D(product_31__N_2324[1]), .SP(w_clk_cpu_enable_711), 
            .CK(w_clk_cpu), .Q(product[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam product_i0_i1.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i26 (.D(\d_result_0[26] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[26])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i26.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i25 (.D(\d_result_0[25] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[25])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i25.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i24 (.D(\d_result_0[24] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[24])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i24.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i23 (.D(\d_result_0[23] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[23])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i23.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i22 (.D(\d_result_0[22] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[22])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i22.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i21 (.D(\d_result_0[21] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[21])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i21.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i20 (.D(\d_result_0[20] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[20])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i20.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i19 (.D(\d_result_0[19] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[19])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i19.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i18 (.D(\d_result_0[18] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[18])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i18.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i17 (.D(\d_result_0[17] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[17])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i17.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i16 (.D(\d_result_0[16] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[16])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i16.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i15 (.D(\d_result_0[15] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[15])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i15.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i14 (.D(\d_result_0[14] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[14])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i14.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i13 (.D(\d_result_0[13] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[13])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i13.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i12 (.D(\d_result_0[12] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[12])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i12.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i11 (.D(\d_result_0[11] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[11])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i11.GSR = "ENABLED";
    FADD2B mult_32u_32u_0_add_5_6 (.A0(mult_32u_32u_0_pp_10_31), .A1(mult_32u_32u_0_pp_10_32), 
           .B0(mult_32u_32u_0_pp_11_31), .B1(mult_32u_32u_0_pp_11_32), .CI(co_mult_32u_32u_0_5_5), 
           .S0(s_mult_32u_32u_0_5_31), .S1(s_mult_32u_32u_0_5_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1P3AX muliplicand_i0_i10 (.D(\d_result_0[10] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[10])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i10.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i9 (.D(\d_result_0[9] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[9])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i9.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i8 (.D(\d_result_0[8] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[8])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i8.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i7 (.D(\d_result_0[7] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[7])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i7.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i6 (.D(\d_result_0[6] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[6])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i6.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i5 (.D(\d_result_0[5] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[5])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i5.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i4 (.D(\d_result_0[4] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i4.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i3 (.D(\d_result_0[3] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i3.GSR = "ENABLED";
    FD1P3AX muliplicand_i0_i2 (.D(\d_result_0[2] ), .SP(w_clk_cpu_enable_984), 
            .CK(w_clk_cpu), .Q(muliplicand[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam muliplicand_i0_i2.GSR = "ENABLED";
    FADD2B mult_32u_32u_0_add_5_5 (.A0(mult_32u_32u_0_pp_10_29), .A1(mult_32u_32u_0_pp_10_30), 
           .B0(mult_32u_32u_0_pp_11_29), .B1(mult_32u_32u_0_pp_11_30), .CI(co_mult_32u_32u_0_5_4), 
           .COUT(co_mult_32u_32u_0_5_5), .S0(s_mult_32u_32u_0_5_29), .S1(s_mult_32u_32u_0_5_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_5_4 (.A0(mult_32u_32u_0_pp_10_27), .A1(mult_32u_32u_0_pp_10_28), 
           .B0(mult_32u_32u_0_pp_11_27), .B1(mult_32u_32u_0_pp_11_28), .CI(co_mult_32u_32u_0_5_3), 
           .COUT(co_mult_32u_32u_0_5_4), .S0(s_mult_32u_32u_0_5_27), .S1(s_mult_32u_32u_0_5_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_5_3 (.A0(mult_32u_32u_0_pp_10_25), .A1(mult_32u_32u_0_pp_10_26), 
           .B0(mult_32u_32u_0_pp_11_25), .B1(mult_32u_32u_0_pp_11_26), .CI(co_mult_32u_32u_0_5_2), 
           .COUT(co_mult_32u_32u_0_5_3), .S0(s_mult_32u_32u_0_5_25), .S1(s_mult_32u_32u_0_5_26)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_6_4 (.A0(mult_32u_32u_0_pp_12_31), .A1(mult_32u_32u_0_pp_12_32), 
           .B0(mult_32u_32u_0_pp_13_31), .B1(mult_32u_32u_0_pp_13_32), .CI(co_mult_32u_32u_0_6_3), 
           .S0(s_mult_32u_32u_0_6_31), .S1(s_mult_32u_32u_0_6_32)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FADD2B mult_32u_32u_0_add_6_3 (.A0(mult_32u_32u_0_pp_12_29), .A1(mult_32u_32u_0_pp_12_30), 
           .B0(mult_32u_32u_0_pp_13_29), .B1(mult_32u_32u_0_pp_13_30), .CI(co_mult_32u_32u_0_6_2), 
           .COUT(co_mult_32u_32u_0_6_3), .S0(s_mult_32u_32u_0_6_29), .S1(s_mult_32u_32u_0_6_30)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1S3AX result_i31 (.D(product[31]), .CK(w_clk_cpu), .Q(multiplier_result_w[31])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i31.GSR = "ENABLED";
    FD1S3AX result_i30 (.D(product[30]), .CK(w_clk_cpu), .Q(multiplier_result_w[30])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i30.GSR = "ENABLED";
    FADD2B mult_32u_32u_0_add_5_2 (.A0(mult_32u_32u_0_pp_10_23), .A1(mult_32u_32u_0_pp_10_24), 
           .B0(mult_32u_32u_0_pp_11_23), .B1(mult_32u_32u_0_pp_11_24), .CI(co_mult_32u_32u_0_5_1), 
           .COUT(co_mult_32u_32u_0_5_2), .S0(s_mult_32u_32u_0_5_23), .S1(s_mult_32u_32u_0_5_24)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1S3AX result_i29 (.D(product[29]), .CK(w_clk_cpu), .Q(multiplier_result_w[29])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i29.GSR = "ENABLED";
    FADD2B mult_32u_32u_0_add_6_2 (.A0(mult_32u_32u_0_pp_12_27), .A1(mult_32u_32u_0_pp_12_28), 
           .B0(mult_32u_32u_0_pp_13_27), .B1(mult_32u_32u_0_pp_13_28), .CI(co_mult_32u_32u_0_6_1), 
           .COUT(co_mult_32u_32u_0_6_2), .S0(s_mult_32u_32u_0_6_27), .S1(s_mult_32u_32u_0_6_28)) /* synthesis syn_instantiated=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(115[27:51])
    FD1S3AX result_i28 (.D(product[28]), .CK(w_clk_cpu), .Q(multiplier_result_w[28])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i28.GSR = "ENABLED";
    FD1S3AX result_i27 (.D(product[27]), .CK(w_clk_cpu), .Q(multiplier_result_w[27])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=1087, LSE_RLINE=1097 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_multiplier.v(108[5] 117[8])
    defparam result_i27.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module lm32_mc_arithmetic
//

module lm32_mc_arithmetic (reg_data_1, w_result, n18863, operand_m, 
            left_shift_result, m_result_sel_shift_m, n1826, n18875, 
            w_clk_cpu, w_clk_cpu_enable_958, n41406, n37259, n41391, 
            load_x, n39970, bypass_data_0, n41417, w_clk_cpu_enable_865, 
            mc_result_x, mc_stall_request_x, GND_net, n21435, n21434, 
            n21433, n21432, n21431, n21430, n21429, n1857, n1856, 
            n1855, n1854, n1853, n41364, n22236, \instruction_d[11] , 
            n41380, n2, n1852, n18869, \instruction_d[12] , n2_adj_50, 
            n1851, \instruction_d[13] , n2_adj_51, \instruction_d[14] , 
            n2_adj_52, sign_extend_immediate, \instruction_d[15] , n36772, 
            \instruction_d[0] , n2_adj_53, \instruction_d[1] , n2_adj_54, 
            \instruction_d[2] , n2_adj_55, \instruction_d[3] , n2_adj_56, 
            \instruction_d[4] , n2_adj_57, \instruction_d[5] , n2_adj_58, 
            \instruction_d[6] , n2_adj_59, \instruction_d[7] , n2_adj_60, 
            \instruction_d[8] , n2_adj_61, \instruction_d[9] , n2_adj_62, 
            \instruction_d[10] , n2_adj_63, divide_by_zero_x, condition_met_m, 
            m_result_sel_compare_m, n41367, raw_x_1, cycles_5__N_2495, 
            csr_read_data_x, adder_result_x, x_result_sel_add_x, \x_result_31__N_616[1] , 
            \x_result_31__N_616[2] , \x_result_31__N_616[3] , \x_result_31__N_616[4] , 
            \x_result_31__N_616[5] , \x_result_31__N_616[6] , \x_result_31__N_616[7] , 
            \x_result_31__N_616[15] , n13, \x_result_31__N_616[16] , \x_result_31__N_616[17] , 
            n41373, n41408, \x_result_31__N_616[18] , \x_result_31__N_616[19] , 
            \x_result_31__N_616[20] , \x_result_31__N_616[21] , \x_result_31__N_616[22] , 
            x_result_sel_csr_x, x_result_sel_sext_x, n41411, direction_m, 
            n41407, pc_f, \x_result_31__N_616[23] , \x_result_31__N_616[24] , 
            \x_result_31__N_616[25] , n42740, n41361, \x_result_31__N_616[26] , 
            \x_result_31__N_616[27] , \x_result_31__N_616[28] , \x_result_31__N_616[0] , 
            \x_result_31__N_616[29] , \x_result_31__N_616[30] , \x_result_31__N_616[31] , 
            w_clk_cpu_enable_984, LM32I_CYC_O, i_cyc_o_N_1759, w_clk_cpu_enable_216, 
            n21414, n37179, \muliplicand[0] , n1285, \muliplicand[7] , 
            \muliplicand[6] , \muliplicand[5] , \muliplicand[4] , \muliplicand[3] , 
            n41345, \muliplicand[2] , \muliplicand[1] , n1844, n1845, 
            n1846, n1847, n38799, n38840, n1791, n1790, n1789, 
            n1788, n1787, n1786, n1785, n1777, n1776, n1775, n1774, 
            n1773, n1772, n1771, n1770, n1769, n1768, n1767, n1766, 
            n1765, n1764, n1792, n1763, n1762, n1843, n1842, n1841, 
            n1840, n1839, n1838, n1837, n1836, n1835) /* synthesis syn_module_defined=1 */ ;
    input [31:0]reg_data_1;
    input [31:0]w_result;
    input n18863;
    input [31:0]operand_m;
    input [31:0]left_shift_result;
    input m_result_sel_shift_m;
    input [31:0]n1826;
    input n18875;
    input w_clk_cpu;
    input w_clk_cpu_enable_958;
    input n41406;
    input n37259;
    input n41391;
    input load_x;
    output n39970;
    input [31:0]bypass_data_0;
    input n41417;
    input w_clk_cpu_enable_865;
    output [31:0]mc_result_x;
    input mc_stall_request_x;
    input GND_net;
    input n21435;
    input n21434;
    input n21433;
    input n21432;
    input n21431;
    input n21430;
    input n21429;
    input n1857;
    input n1856;
    input n1855;
    input n1854;
    input n1853;
    input n41364;
    input n22236;
    input \instruction_d[11] ;
    input n41380;
    output n2;
    input n1852;
    input n18869;
    input \instruction_d[12] ;
    output n2_adj_50;
    input n1851;
    input \instruction_d[13] ;
    output n2_adj_51;
    input \instruction_d[14] ;
    output n2_adj_52;
    input sign_extend_immediate;
    input \instruction_d[15] ;
    output n36772;
    input \instruction_d[0] ;
    output n2_adj_53;
    input \instruction_d[1] ;
    output n2_adj_54;
    input \instruction_d[2] ;
    output n2_adj_55;
    input \instruction_d[3] ;
    output n2_adj_56;
    input \instruction_d[4] ;
    output n2_adj_57;
    input \instruction_d[5] ;
    output n2_adj_58;
    input \instruction_d[6] ;
    output n2_adj_59;
    input \instruction_d[7] ;
    output n2_adj_60;
    input \instruction_d[8] ;
    output n2_adj_61;
    input \instruction_d[9] ;
    output n2_adj_62;
    input \instruction_d[10] ;
    output n2_adj_63;
    output divide_by_zero_x;
    input condition_met_m;
    input m_result_sel_compare_m;
    input n41367;
    input raw_x_1;
    output cycles_5__N_2495;
    input [31:0]csr_read_data_x;
    input [31:0]adder_result_x;
    input x_result_sel_add_x;
    output \x_result_31__N_616[1] ;
    output \x_result_31__N_616[2] ;
    output \x_result_31__N_616[3] ;
    output \x_result_31__N_616[4] ;
    output \x_result_31__N_616[5] ;
    output \x_result_31__N_616[6] ;
    output \x_result_31__N_616[7] ;
    output \x_result_31__N_616[15] ;
    output n13;
    output \x_result_31__N_616[16] ;
    output \x_result_31__N_616[17] ;
    input n41373;
    input n41408;
    output \x_result_31__N_616[18] ;
    output \x_result_31__N_616[19] ;
    output \x_result_31__N_616[20] ;
    output \x_result_31__N_616[21] ;
    output \x_result_31__N_616[22] ;
    input x_result_sel_csr_x;
    input x_result_sel_sext_x;
    input n41411;
    input direction_m;
    input n41407;
    input [31:2]pc_f;
    output \x_result_31__N_616[23] ;
    output \x_result_31__N_616[24] ;
    output \x_result_31__N_616[25] ;
    input n42740;
    input n41361;
    output \x_result_31__N_616[26] ;
    output \x_result_31__N_616[27] ;
    output \x_result_31__N_616[28] ;
    output \x_result_31__N_616[0] ;
    output \x_result_31__N_616[29] ;
    output \x_result_31__N_616[30] ;
    output \x_result_31__N_616[31] ;
    input w_clk_cpu_enable_984;
    input LM32I_CYC_O;
    input i_cyc_o_N_1759;
    output w_clk_cpu_enable_216;
    input n21414;
    output n37179;
    input \muliplicand[0] ;
    input n1285;
    input \muliplicand[7] ;
    input \muliplicand[6] ;
    input \muliplicand[5] ;
    input \muliplicand[4] ;
    input \muliplicand[3] ;
    input n41345;
    input \muliplicand[2] ;
    input \muliplicand[1] ;
    input n1844;
    input n1845;
    input n1846;
    input n1847;
    input n38799;
    input n38840;
    input n1791;
    input n1790;
    input n1789;
    input n1788;
    input n1787;
    input n1786;
    input n1785;
    input n1777;
    input n1776;
    input n1775;
    input n1774;
    input n1773;
    input n1772;
    input n1771;
    input n1770;
    input n1769;
    input n1768;
    input n1767;
    input n1766;
    input n1765;
    input n1764;
    input n1792;
    input n1763;
    input n1762;
    input n1843;
    input n1842;
    input n1841;
    input n1840;
    input n1839;
    input n1838;
    input n1837;
    input n1836;
    input n1835;
    
    wire w_clk_cpu /* synthesis SET_AS_NETWORK=w_clk_cpu, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(22[6:15])
    wire [31:0]n1562;
    wire [31:0]n1595;
    
    wire n41301;
    wire [31:0]n1900;
    wire [31:0]n1793;
    wire [31:0]b;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(134[22:23])
    
    wire n22517;
    wire [31:0]n1976;
    
    wire n40484, n40477, n40478;
    wire [31:0]a;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(133[22:23])
    wire [31:0]n18884;
    
    wire n40476;
    wire [31:0]n1461;
    
    wire n40483, n40482, n36638;
    wire [31:0]p;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(132[22:23])
    wire [32:0]t;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(136[13:14])
    
    wire n36639;
    wire [31:0]n1727;
    
    wire n18873;
    wire [31:0]n1862;
    
    wire n36637, n36636;
    wire [2:0]state;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(139[26:31])
    wire [31:0]n1826_c;
    
    wire n41317, n41316, n41318, n41314, n41313, n41315, n41306, 
        n41305, n41307;
    wire [5:0]cycles;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(140[11:17])
    wire [5:0]n29;
    
    wire n41303, n41302, n41304, cycles_5__N_2497, n23934, n41300, 
        n41299, divide_by_zero_x_N_2647;
    wire [31:0]n19597;
    wire [31:0]n1628;
    wire [31:0]n18918;
    
    wire n4, n9, n18879, n23940, n23938;
    wire [5:0]n37;
    
    wire n16, n24948, divide_by_zero_x_N_2651, n10, n18877;
    wire [31:0]n1936;
    
    wire n24658, n39272, n4_adj_3775, n39274, n39270, n39244, n39128, 
        n39108, n39266, n39236, n39104, n39240, n39118, n39232, 
        n39094, n36661, n36660, n36659, n36651, n36650, n36649, 
        n36648, n36647, n36646, n36645, n36644, n36643, n36642, 
        n36641, n36640;
    
    LUT4 mux_675_i18_3_lut (.A(reg_data_1[17]), .B(w_result[17]), .C(n18863), 
         .Z(n1562[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i18_3_lut.init = 16'hcaca;
    LUT4 mux_676_i17_3_lut (.A(operand_m[16]), .B(left_shift_result[15]), 
         .C(m_result_sel_shift_m), .Z(n1595[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i17_3_lut.init = 16'hcaca;
    LUT4 i37768_3_lut (.A(n41301), .B(n1826[10]), .C(n18875), .Z(n1900[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37768_3_lut.init = 16'hcaca;
    LUT4 mux_675_i17_3_lut (.A(reg_data_1[16]), .B(w_result[16]), .C(n18863), 
         .Z(n1562[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i17_3_lut.init = 16'hcaca;
    PFUMX mux_693_i25 (.BLUT(n1793[24]), .ALUT(n1826[24]), .C0(n18875), 
          .Z(n1900[24]));
    LUT4 mux_676_i16_3_lut (.A(operand_m[15]), .B(left_shift_result[16]), 
         .C(m_result_sel_shift_m), .Z(n1595[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i16_3_lut.init = 16'hcaca;
    LUT4 mux_675_i16_3_lut (.A(reg_data_1[15]), .B(w_result[15]), .C(n18863), 
         .Z(n1562[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i16_3_lut.init = 16'hcaca;
    FD1P3IX b__i20 (.D(n1976[20]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[20])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i20.GSR = "ENABLED";
    LUT4 i37770_3_lut (.A(n40484), .B(n1826[9]), .C(n18875), .Z(n1900[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37770_3_lut.init = 16'hcaca;
    FD1P3IX b__i5 (.D(n1976[5]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[5])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i5.GSR = "ENABLED";
    FD1P3IX b__i31 (.D(n1976[31]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[31])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i31.GSR = "ENABLED";
    PFUMX mux_693_i26 (.BLUT(n1793[25]), .ALUT(n1826[25]), .C0(n18875), 
          .Z(n1900[25]));
    FD1P3IX b__i19 (.D(n1976[19]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[19])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i19.GSR = "ENABLED";
    FD1P3IX b__i4 (.D(n1976[4]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i4.GSR = "ENABLED";
    FD1P3IX b__i30 (.D(n1976[30]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[30])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i30.GSR = "ENABLED";
    LUT4 reg_data_1_8__bdd_3_lut_39255 (.A(reg_data_1[8]), .B(w_result[8]), 
         .C(n18863), .Z(n40477)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam reg_data_1_8__bdd_3_lut_39255.init = 16'hcaca;
    FD1P3IX b__i18 (.D(n1976[18]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[18])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i18.GSR = "ENABLED";
    FD1P3IX b__i3 (.D(n1976[3]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i3.GSR = "ENABLED";
    LUT4 i37888_4_lut (.A(n41406), .B(n37259), .C(n41391), .D(load_x), 
         .Z(n39970)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2265[34:53])
    defparam i37888_4_lut.init = 16'h1333;
    LUT4 i37772_3_lut (.A(n40478), .B(n1826[8]), .C(n18875), .Z(n1900[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37772_3_lut.init = 16'hcaca;
    LUT4 mux_17581_i2_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[1]), 
         .C(a[0]), .D(n41417), .Z(n18884[1])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i2_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 reg_data_1_8__bdd_3_lut_38122 (.A(operand_m[8]), .B(m_result_sel_shift_m), 
         .C(left_shift_result[23]), .Z(n40476)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam reg_data_1_8__bdd_3_lut_38122.init = 16'he2e2;
    FD1P3IX a_i0_i1 (.D(n18884[1]), .SP(w_clk_cpu_enable_865), .CD(n22517), 
            .CK(w_clk_cpu), .Q(a[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i1.GSR = "ENABLED";
    FD1P3IX b__i17 (.D(n1976[17]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[17])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i17.GSR = "ENABLED";
    FD1P3AX result_x_i0_i3 (.D(n1461[3]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i3.GSR = "ENABLED";
    FD1P3AX result_x_i0_i2 (.D(n1461[2]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i2.GSR = "ENABLED";
    FD1P3IX b__i2 (.D(n1976[2]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i2.GSR = "ENABLED";
    PFUMX mux_693_i27 (.BLUT(n1793[26]), .ALUT(n1826[26]), .C0(n18875), 
          .Z(n1900[26]));
    LUT4 reg_data_1_9__bdd_3_lut_39263 (.A(reg_data_1[9]), .B(w_result[9]), 
         .C(n18863), .Z(n40483)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam reg_data_1_9__bdd_3_lut_39263.init = 16'hcaca;
    FD1P3IX b__i16 (.D(n1976[16]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[16])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i16.GSR = "ENABLED";
    FD1P3IX b__i1 (.D(n1976[1]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i1.GSR = "ENABLED";
    PFUMX mux_693_i28 (.BLUT(n1793[27]), .ALUT(n1826[27]), .C0(n18875), 
          .Z(n1900[27]));
    FD1P3IX b__i0 (.D(n1976[0]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i0.GSR = "ENABLED";
    LUT4 reg_data_1_9__bdd_3_lut_38127 (.A(operand_m[9]), .B(m_result_sel_shift_m), 
         .C(left_shift_result[22]), .Z(n40482)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam reg_data_1_9__bdd_3_lut_38127.init = 16'he2e2;
    PFUMX mux_693_i29 (.BLUT(n1793[28]), .ALUT(n1826[28]), .C0(n18875), 
          .Z(n1900[28]));
    FD1P3AX result_x_i0_i1 (.D(n1461[1]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i1.GSR = "ENABLED";
    PFUMX mux_693_i30 (.BLUT(n1793[29]), .ALUT(n1826[29]), .C0(n18875), 
          .Z(n1900[29]));
    FD1P3IX b__i29 (.D(n1976[29]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[29])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i29.GSR = "ENABLED";
    PFUMX mux_693_i31 (.BLUT(n1793[30]), .ALUT(n1826[30]), .C0(n18875), 
          .Z(n1900[30]));
    CCU2D p_30__I_0_add_2_7 (.A0(p[4]), .B0(b[5]), .C0(GND_net), .D0(GND_net), 
          .A1(p[5]), .B1(b[6]), .C1(GND_net), .D1(GND_net), .CIN(n36638), 
          .COUT(n36639), .S0(t[5]), .S1(t[6]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam p_30__I_0_add_2_7.INIT0 = 16'h5999;
    defparam p_30__I_0_add_2_7.INIT1 = 16'h5999;
    defparam p_30__I_0_add_2_7.INJECT1_0 = "NO";
    defparam p_30__I_0_add_2_7.INJECT1_1 = "NO";
    PFUMX mux_693_i32 (.BLUT(n1793[31]), .ALUT(n1826[31]), .C0(n18875), 
          .Z(n1900[31]));
    PFUMX mux_687_i9 (.BLUT(n21435), .ALUT(n1727[8]), .C0(n18873), .Z(n1862[8]));
    PFUMX mux_687_i10 (.BLUT(n21434), .ALUT(n1727[9]), .C0(n18873), .Z(n1862[9]));
    CCU2D p_30__I_0_add_2_5 (.A0(p[2]), .B0(b[3]), .C0(GND_net), .D0(GND_net), 
          .A1(p[3]), .B1(b[4]), .C1(GND_net), .D1(GND_net), .CIN(n36637), 
          .COUT(n36638), .S0(t[3]), .S1(t[4]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam p_30__I_0_add_2_5.INIT0 = 16'h5999;
    defparam p_30__I_0_add_2_5.INIT1 = 16'h5999;
    defparam p_30__I_0_add_2_5.INJECT1_0 = "NO";
    defparam p_30__I_0_add_2_5.INJECT1_1 = "NO";
    FD1P3IX b__i15 (.D(n1976[15]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[15])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i15.GSR = "ENABLED";
    PFUMX mux_687_i11 (.BLUT(n21433), .ALUT(n1727[10]), .C0(n18873), .Z(n1862[10]));
    PFUMX mux_687_i12 (.BLUT(n21432), .ALUT(n1727[11]), .C0(n18873), .Z(n1862[11]));
    PFUMX mux_687_i13 (.BLUT(n21431), .ALUT(n1727[12]), .C0(n18873), .Z(n1862[12]));
    CCU2D p_30__I_0_add_2_3 (.A0(p[0]), .B0(b[1]), .C0(GND_net), .D0(GND_net), 
          .A1(p[1]), .B1(b[2]), .C1(GND_net), .D1(GND_net), .CIN(n36636), 
          .COUT(n36637), .S0(t[1]), .S1(t[2]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam p_30__I_0_add_2_3.INIT0 = 16'h5999;
    defparam p_30__I_0_add_2_3.INIT1 = 16'h5999;
    defparam p_30__I_0_add_2_3.INJECT1_0 = "NO";
    defparam p_30__I_0_add_2_3.INJECT1_1 = "NO";
    PFUMX mux_687_i14 (.BLUT(n21430), .ALUT(n1727[13]), .C0(n18873), .Z(n1862[13]));
    PFUMX mux_687_i15 (.BLUT(n21429), .ALUT(n1727[14]), .C0(n18873), .Z(n1862[14]));
    LUT4 mux_670_i2_3_lut (.A(p[1]), .B(a[1]), .C(state[0]), .Z(n1461[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i2_3_lut.init = 16'hcaca;
    PFUMX mux_693_i1 (.BLUT(n1793[0]), .ALUT(n1826_c[0]), .C0(n18875), 
          .Z(n1900[0]));
    PFUMX mux_693_i2 (.BLUT(n1793[1]), .ALUT(n1857), .C0(n18875), .Z(n1900[1]));
    CCU2D p_30__I_0_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(a[31]), .B1(b[0]), .C1(GND_net), .D1(GND_net), 
          .COUT(n36636), .S1(t[0]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam p_30__I_0_add_2_1.INIT0 = 16'h0000;
    defparam p_30__I_0_add_2_1.INIT1 = 16'h5999;
    defparam p_30__I_0_add_2_1.INJECT1_0 = "NO";
    defparam p_30__I_0_add_2_1.INJECT1_1 = "NO";
    PFUMX mux_693_i3 (.BLUT(n1793[2]), .ALUT(n1856), .C0(n18875), .Z(n1900[2]));
    PFUMX mux_693_i4 (.BLUT(n1793[3]), .ALUT(n1855), .C0(n18875), .Z(n1900[3]));
    PFUMX mux_693_i5 (.BLUT(n1793[4]), .ALUT(n1854), .C0(n18875), .Z(n1900[4]));
    PFUMX mux_693_i6 (.BLUT(n1793[5]), .ALUT(n1853), .C0(n18875), .Z(n1900[5]));
    LUT4 i28879_4_lut_4_lut (.A(n41364), .B(n22236), .C(\instruction_d[11] ), 
         .D(n41380), .Z(n2)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;
    defparam i28879_4_lut_4_lut.init = 16'h5140;
    PFUMX mux_693_i7 (.BLUT(n1793[6]), .ALUT(n1852), .C0(n18875), .Z(n1900[6]));
    PFUMX i38545 (.BLUT(n41317), .ALUT(n41316), .C0(n18869), .Z(n41318));
    LUT4 mux_17581_i32_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[31]), 
         .C(a[30]), .D(n41417), .Z(n18884[31])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i32_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i28880_4_lut_4_lut (.A(n41364), .B(n22236), .C(\instruction_d[12] ), 
         .D(n41380), .Z(n2_adj_50)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;
    defparam i28880_4_lut_4_lut.init = 16'h5140;
    LUT4 mux_17581_i31_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[30]), 
         .C(a[29]), .D(n41417), .Z(n18884[30])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i31_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 mux_17581_i30_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[29]), 
         .C(a[28]), .D(n41417), .Z(n18884[29])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i30_3_lut_4_lut_4_lut.init = 16'hf0d8;
    PFUMX mux_693_i8 (.BLUT(n1793[7]), .ALUT(n1851), .C0(n18875), .Z(n1900[7]));
    LUT4 i28891_4_lut_4_lut (.A(n41364), .B(n22236), .C(\instruction_d[13] ), 
         .D(n41380), .Z(n2_adj_51)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;
    defparam i28891_4_lut_4_lut.init = 16'h5140;
    PFUMX i38542 (.BLUT(n41314), .ALUT(n41313), .C0(n18869), .Z(n41315));
    LUT4 i28899_4_lut_4_lut (.A(n41364), .B(n22236), .C(\instruction_d[14] ), 
         .D(n41380), .Z(n2_adj_52)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;
    defparam i28899_4_lut_4_lut.init = 16'h5140;
    LUT4 i2_4_lut_4_lut (.A(n41364), .B(sign_extend_immediate), .C(n22236), 
         .D(\instruction_d[15] ), .Z(n36772)) /* synthesis lut_function=(!(A+!(B (D)+!B (C (D))))) */ ;
    defparam i2_4_lut_4_lut.init = 16'h5400;
    LUT4 i29640_4_lut_4_lut (.A(n41364), .B(n22236), .C(\instruction_d[0] ), 
         .D(n41380), .Z(n2_adj_53)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;
    defparam i29640_4_lut_4_lut.init = 16'h5140;
    LUT4 i29647_4_lut_4_lut (.A(n41364), .B(n22236), .C(\instruction_d[1] ), 
         .D(n41380), .Z(n2_adj_54)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;
    defparam i29647_4_lut_4_lut.init = 16'h5140;
    LUT4 mux_17581_i29_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[28]), 
         .C(a[27]), .D(n41417), .Z(n18884[28])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i29_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 mux_17581_i28_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[27]), 
         .C(a[26]), .D(n41417), .Z(n18884[27])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i28_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i29660_4_lut_4_lut (.A(n41364), .B(n22236), .C(\instruction_d[2] ), 
         .D(n41380), .Z(n2_adj_55)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;
    defparam i29660_4_lut_4_lut.init = 16'h5140;
    LUT4 i29668_4_lut_4_lut (.A(n41364), .B(n22236), .C(\instruction_d[3] ), 
         .D(n41380), .Z(n2_adj_56)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;
    defparam i29668_4_lut_4_lut.init = 16'h5140;
    LUT4 i29680_4_lut_4_lut (.A(n41364), .B(n22236), .C(\instruction_d[4] ), 
         .D(n41380), .Z(n2_adj_57)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;
    defparam i29680_4_lut_4_lut.init = 16'h5140;
    LUT4 i29688_4_lut_4_lut (.A(n41364), .B(n22236), .C(\instruction_d[5] ), 
         .D(n41380), .Z(n2_adj_58)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;
    defparam i29688_4_lut_4_lut.init = 16'h5140;
    LUT4 i29697_4_lut_4_lut (.A(n41364), .B(n22236), .C(\instruction_d[6] ), 
         .D(n41380), .Z(n2_adj_59)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;
    defparam i29697_4_lut_4_lut.init = 16'h5140;
    LUT4 i29704_4_lut_4_lut (.A(n41364), .B(n22236), .C(\instruction_d[7] ), 
         .D(n41380), .Z(n2_adj_60)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;
    defparam i29704_4_lut_4_lut.init = 16'h5140;
    LUT4 i29714_4_lut_4_lut (.A(n41364), .B(n22236), .C(\instruction_d[8] ), 
         .D(n41380), .Z(n2_adj_61)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;
    defparam i29714_4_lut_4_lut.init = 16'h5140;
    LUT4 mux_17581_i27_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[26]), 
         .C(a[25]), .D(n41417), .Z(n18884[26])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i27_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 mux_17581_i26_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[25]), 
         .C(a[24]), .D(n41417), .Z(n18884[25])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i26_3_lut_4_lut_4_lut.init = 16'hf0d8;
    PFUMX i38536 (.BLUT(n41306), .ALUT(n41305), .C0(n18869), .Z(n41307));
    LUT4 i29722_4_lut_4_lut (.A(n41364), .B(n22236), .C(\instruction_d[9] ), 
         .D(n41380), .Z(n2_adj_62)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;
    defparam i29722_4_lut_4_lut.init = 16'h5140;
    LUT4 i28827_4_lut_4_lut (.A(n41364), .B(n22236), .C(\instruction_d[10] ), 
         .D(n41380), .Z(n2_adj_63)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;
    defparam i28827_4_lut_4_lut.init = 16'h5140;
    FD1P3IX cycles_19669__i1 (.D(n29[1]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(cycles[1])) /* synthesis syn_use_carry_chain=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(250[26:39])
    defparam cycles_19669__i1.GSR = "ENABLED";
    LUT4 mux_17581_i25_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[24]), 
         .C(a[23]), .D(n41417), .Z(n18884[24])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i25_3_lut_4_lut_4_lut.init = 16'hf0d8;
    FD1P3IX b__i28 (.D(n1976[28]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[28])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i28.GSR = "ENABLED";
    FD1P3IX b__i14 (.D(n1976[14]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[14])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i14.GSR = "ENABLED";
    FD1P3IX b__i27 (.D(n1976[27]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[27])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i27.GSR = "ENABLED";
    PFUMX i38533 (.BLUT(n41303), .ALUT(n41302), .C0(n18869), .Z(n41304));
    FD1P3IX b__i13 (.D(n1976[13]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[13])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i13.GSR = "ENABLED";
    FD1S3AX state_FSM_i1 (.D(n23934), .CK(w_clk_cpu), .Q(cycles_5__N_2497));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam state_FSM_i1.GSR = "ENABLED";
    LUT4 mux_17581_i24_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[23]), 
         .C(a[22]), .D(n41417), .Z(n18884[23])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i24_3_lut_4_lut_4_lut.init = 16'hf0d8;
    PFUMX i38530 (.BLUT(n41300), .ALUT(n41299), .C0(n18869), .Z(n41301));
    LUT4 mux_17581_i23_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[22]), 
         .C(a[21]), .D(n41417), .Z(n18884[22])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i23_3_lut_4_lut_4_lut.init = 16'hf0d8;
    FD1P3IX cycles_19669__i2 (.D(n29[2]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(cycles[2])) /* synthesis syn_use_carry_chain=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(250[26:39])
    defparam cycles_19669__i2.GSR = "ENABLED";
    FD1P3IX b__i26 (.D(n1976[26]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[26])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i26.GSR = "ENABLED";
    FD1P3IX b__i12 (.D(n1976[12]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[12])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i12.GSR = "ENABLED";
    FD1P3IX b__i25 (.D(n1976[25]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[25])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i25.GSR = "ENABLED";
    FD1P3IX b__i11 (.D(n1976[11]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[11])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i11.GSR = "ENABLED";
    FD1P3IX cycles_19669__i3 (.D(n29[3]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(cycles[3])) /* synthesis syn_use_carry_chain=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(250[26:39])
    defparam cycles_19669__i3.GSR = "ENABLED";
    FD1P3IX cycles_19669__i4 (.D(n29[4]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(cycles[4])) /* synthesis syn_use_carry_chain=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(250[26:39])
    defparam cycles_19669__i4.GSR = "ENABLED";
    LUT4 mux_17581_i22_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[21]), 
         .C(a[20]), .D(n41417), .Z(n18884[21])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i22_3_lut_4_lut_4_lut.init = 16'hf0d8;
    FD1P3AX result_x_i0_i0 (.D(n1461[0]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i0.GSR = "ENABLED";
    FD1S3AX divide_by_zero_x_58 (.D(divide_by_zero_x_N_2647), .CK(w_clk_cpu), 
            .Q(divide_by_zero_x)) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam divide_by_zero_x_58.GSR = "ENABLED";
    LUT4 mux_17581_i21_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[20]), 
         .C(a[19]), .D(n41417), .Z(n18884[20])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i21_3_lut_4_lut_4_lut.init = 16'hf0d8;
    FD1P3IX b__i10 (.D(n1976[10]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[10])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i10.GSR = "ENABLED";
    FD1P3IX cycles_19669__i0 (.D(n29[0]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(cycles[0])) /* synthesis syn_use_carry_chain=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(250[26:39])
    defparam cycles_19669__i0.GSR = "ENABLED";
    LUT4 mux_17581_i20_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[19]), 
         .C(a[18]), .D(n41417), .Z(n18884[19])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i20_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 mux_17581_i19_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[18]), 
         .C(a[17]), .D(n41417), .Z(n18884[18])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i19_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 mux_17581_i18_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[17]), 
         .C(a[16]), .D(n41417), .Z(n18884[17])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i18_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 mux_17581_i17_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[16]), 
         .C(a[15]), .D(n41417), .Z(n18884[16])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i17_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 mux_17581_i1_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[0]), 
         .C(t[32]), .D(n41417), .Z(n18884[0])) /* synthesis lut_function=(!(A (B (C (D))+!B (C+!(D)))+!A (C))) */ ;
    defparam mux_17581_i1_3_lut_4_lut_4_lut.init = 16'h0f8d;
    LUT4 mux_18230_i32_3_lut (.A(t[31]), .B(p[30]), .C(t[32]), .Z(n19597[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i32_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i31_3_lut (.A(t[30]), .B(p[29]), .C(t[32]), .Z(n19597[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i31_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i30_3_lut (.A(t[29]), .B(p[28]), .C(t[32]), .Z(n19597[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i30_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i29_3_lut (.A(t[28]), .B(p[27]), .C(t[32]), .Z(n19597[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i29_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i28_3_lut (.A(t[27]), .B(p[26]), .C(t[32]), .Z(n19597[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i28_3_lut.init = 16'hcaca;
    FD1P3IX b__i24 (.D(n1976[24]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[24])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i24.GSR = "ENABLED";
    FD1P3IX b__i9 (.D(n1976[9]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[9])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i9.GSR = "ENABLED";
    LUT4 mux_17581_i16_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[15]), 
         .C(a[14]), .D(n41417), .Z(n18884[15])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i16_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 mux_17581_i15_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[14]), 
         .C(a[13]), .D(n41417), .Z(n18884[14])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i15_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 mux_17581_i14_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[13]), 
         .C(a[12]), .D(n41417), .Z(n18884[13])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i14_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 mux_18230_i27_3_lut (.A(t[26]), .B(p[25]), .C(t[32]), .Z(n19597[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i27_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i26_3_lut (.A(t[25]), .B(p[24]), .C(t[32]), .Z(n19597[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i26_3_lut.init = 16'hcaca;
    LUT4 mux_677_i1_3_lut (.A(left_shift_result[0]), .B(condition_met_m), 
         .C(m_result_sel_compare_m), .Z(n1628[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_677_i1_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i25_3_lut (.A(t[24]), .B(p[23]), .C(t[32]), .Z(n19597[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i25_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i24_3_lut (.A(t[23]), .B(p[22]), .C(t[32]), .Z(n19597[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i24_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i23_3_lut (.A(t[22]), .B(p[21]), .C(t[32]), .Z(n19597[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i23_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i22_3_lut (.A(t[21]), .B(p[20]), .C(t[32]), .Z(n19597[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i22_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i1_3_lut (.A(t[0]), .B(a[31]), .C(t[32]), .Z(n19597[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i1_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i21_3_lut (.A(t[20]), .B(p[19]), .C(t[32]), .Z(n19597[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i21_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i20_3_lut (.A(t[19]), .B(p[18]), .C(t[32]), .Z(n19597[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i20_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i19_3_lut (.A(t[18]), .B(p[17]), .C(t[32]), .Z(n19597[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i19_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i18_3_lut (.A(t[17]), .B(p[16]), .C(t[32]), .Z(n19597[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i18_3_lut.init = 16'hcaca;
    FD1P3AX a_i0_i31 (.D(n18918[31]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[31])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i31.GSR = "ENABLED";
    LUT4 mux_18230_i17_3_lut (.A(t[16]), .B(p[15]), .C(t[32]), .Z(n19597[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i17_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i16_3_lut (.A(t[15]), .B(p[14]), .C(t[32]), .Z(n19597[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i16_3_lut.init = 16'hcaca;
    FD1P3AX a_i0_i30 (.D(n18918[30]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[30])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i30.GSR = "ENABLED";
    FD1P3IX p__i0 (.D(n19597[0]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i0.GSR = "ENABLED";
    FD1P3AX a_i0_i29 (.D(n18918[29]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[29])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i29.GSR = "ENABLED";
    LUT4 mux_18230_i15_3_lut (.A(t[14]), .B(p[13]), .C(t[32]), .Z(n19597[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i15_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i14_3_lut (.A(t[13]), .B(p[12]), .C(t[32]), .Z(n19597[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i14_3_lut.init = 16'hcaca;
    FD1P3AX a_i0_i28 (.D(n18918[28]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[28])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i28.GSR = "ENABLED";
    LUT4 mux_17581_i13_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[12]), 
         .C(a[11]), .D(n41417), .Z(n18884[12])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i13_3_lut_4_lut_4_lut.init = 16'hf0d8;
    FD1P3AX a_i0_i27 (.D(n18918[27]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[27])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i27.GSR = "ENABLED";
    LUT4 mux_18230_i13_3_lut (.A(t[12]), .B(p[11]), .C(t[32]), .Z(n19597[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i13_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i12_3_lut (.A(t[11]), .B(p[10]), .C(t[32]), .Z(n19597[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i12_3_lut.init = 16'hcaca;
    LUT4 i37689_3_lut (.A(n1562[23]), .B(n1595[23]), .C(n18869), .Z(n1793[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37689_3_lut.init = 16'hcaca;
    LUT4 i37691_3_lut (.A(n1562[22]), .B(n1595[22]), .C(n18869), .Z(n1793[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37691_3_lut.init = 16'hcaca;
    FD1P3AX a_i0_i26 (.D(n18918[26]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[26])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i26.GSR = "ENABLED";
    LUT4 i37693_3_lut (.A(n1562[21]), .B(n1595[21]), .C(n18869), .Z(n1793[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37693_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut (.A(n41367), .B(n4), .C(raw_x_1), .D(n9), .Z(n18879)) /* synthesis lut_function=(A (B (C (D)))+!A (B)) */ ;
    defparam i2_4_lut.init = 16'hc444;
    FD1P3AX a_i0_i25 (.D(n18918[25]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[25])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i25.GSR = "ENABLED";
    FD1P3AX a_i0_i24 (.D(n18918[24]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[24])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i24.GSR = "ENABLED";
    LUT4 mux_18230_i11_3_lut (.A(t[10]), .B(p[9]), .C(t[32]), .Z(n19597[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i11_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i10_3_lut (.A(t[9]), .B(p[8]), .C(t[32]), .Z(n19597[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i10_3_lut.init = 16'hcaca;
    LUT4 mux_17581_i12_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[11]), 
         .C(a[10]), .D(n41417), .Z(n18884[11])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i12_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 i37695_3_lut (.A(n1562[20]), .B(n1595[20]), .C(n18869), .Z(n1793[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37695_3_lut.init = 16'hcaca;
    FD1P3AX a_i0_i23 (.D(n18918[23]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[23])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i23.GSR = "ENABLED";
    LUT4 mux_17581_i11_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[10]), 
         .C(a[9]), .D(n41417), .Z(n18884[10])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i11_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 mux_18230_i9_3_lut (.A(t[8]), .B(p[7]), .C(t[32]), .Z(n19597[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i9_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i8_3_lut (.A(t[7]), .B(p[6]), .C(t[32]), .Z(n19597[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i8_3_lut.init = 16'hcaca;
    LUT4 mux_670_i32_3_lut (.A(p[31]), .B(a[31]), .C(state[0]), .Z(n1461[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i32_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i7_3_lut (.A(t[6]), .B(p[5]), .C(t[32]), .Z(n19597[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i7_3_lut.init = 16'hcaca;
    FD1P3AX a_i0_i22 (.D(n18918[22]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[22])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i22.GSR = "ENABLED";
    FD1P3AX a_i0_i21 (.D(n18918[21]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[21])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i21.GSR = "ENABLED";
    LUT4 mux_18230_i6_3_lut (.A(t[5]), .B(p[4]), .C(t[32]), .Z(n19597[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i6_3_lut.init = 16'hcaca;
    LUT4 i37697_3_lut (.A(n1562[19]), .B(n1595[19]), .C(n18869), .Z(n1793[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37697_3_lut.init = 16'hcaca;
    FD1P3AX a_i0_i20 (.D(n18918[20]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[20])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i20.GSR = "ENABLED";
    FD1P3AX a_i0_i19 (.D(n18918[19]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[19])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i19.GSR = "ENABLED";
    LUT4 mux_670_i31_3_lut (.A(p[30]), .B(a[30]), .C(state[0]), .Z(n1461[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i31_3_lut.init = 16'hcaca;
    LUT4 mux_670_i30_3_lut (.A(p[29]), .B(a[29]), .C(state[0]), .Z(n1461[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i30_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i5_3_lut (.A(t[4]), .B(p[3]), .C(t[32]), .Z(n19597[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i5_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i4_3_lut (.A(t[3]), .B(p[2]), .C(t[32]), .Z(n19597[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i4_3_lut.init = 16'hcaca;
    LUT4 mux_17581_i10_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[9]), 
         .C(a[8]), .D(n41417), .Z(n18884[9])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i10_3_lut_4_lut_4_lut.init = 16'hf0d8;
    FD1S3AY state_FSM_i3 (.D(n23940), .CK(w_clk_cpu), .Q(cycles_5__N_2495));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam state_FSM_i3.GSR = "ENABLED";
    LUT4 i37699_3_lut (.A(n1562[18]), .B(n1595[18]), .C(n18869), .Z(n1793[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37699_3_lut.init = 16'hcaca;
    FD1P3AX a_i0_i18 (.D(n18918[18]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[18])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i18.GSR = "ENABLED";
    LUT4 mux_670_i29_3_lut (.A(p[28]), .B(a[28]), .C(state[0]), .Z(n1461[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i29_3_lut.init = 16'hcaca;
    LUT4 mux_17581_i9_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[8]), 
         .C(a[7]), .D(n41417), .Z(n18884[8])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i9_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 mux_670_i28_3_lut (.A(p[27]), .B(a[27]), .C(state[0]), .Z(n1461[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i28_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i3_3_lut (.A(t[2]), .B(p[1]), .C(t[32]), .Z(n19597[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i3_3_lut.init = 16'hcaca;
    LUT4 mux_18230_i2_3_lut (.A(t[1]), .B(p[0]), .C(t[32]), .Z(n19597[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_18230_i2_3_lut.init = 16'hcaca;
    LUT4 mux_680_i2_3_lut (.A(csr_read_data_x[1]), .B(adder_result_x[1]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[1] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i2_3_lut.init = 16'hcaca;
    LUT4 mux_680_i3_3_lut (.A(csr_read_data_x[2]), .B(adder_result_x[2]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[2] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i3_3_lut.init = 16'hcaca;
    FD1S3AX state_FSM_i2 (.D(n23938), .CK(w_clk_cpu), .Q(state[0]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam state_FSM_i2.GSR = "ENABLED";
    LUT4 i37701_3_lut (.A(n1562[17]), .B(n1595[17]), .C(n18869), .Z(n1793[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37701_3_lut.init = 16'hcaca;
    FD1P3AX a_i0_i17 (.D(n18918[17]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[17])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i17.GSR = "ENABLED";
    LUT4 mux_670_i27_3_lut (.A(p[26]), .B(a[26]), .C(state[0]), .Z(n1461[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i27_3_lut.init = 16'hcaca;
    LUT4 mux_670_i26_3_lut (.A(p[25]), .B(a[25]), .C(state[0]), .Z(n1461[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i26_3_lut.init = 16'hcaca;
    LUT4 mux_680_i4_3_lut (.A(csr_read_data_x[3]), .B(adder_result_x[3]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[3] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i4_3_lut.init = 16'hcaca;
    LUT4 mux_680_i5_3_lut (.A(csr_read_data_x[4]), .B(adder_result_x[4]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[4] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i5_3_lut.init = 16'hcaca;
    LUT4 mux_680_i6_3_lut (.A(csr_read_data_x[5]), .B(adder_result_x[5]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[5] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i6_3_lut.init = 16'hcaca;
    FD1P3AX a_i0_i16 (.D(n18918[16]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[16])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i16.GSR = "ENABLED";
    FD1P3IX a_i0_i0 (.D(n18884[0]), .SP(w_clk_cpu_enable_865), .CD(n22517), 
            .CK(w_clk_cpu), .Q(a[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i0.GSR = "ENABLED";
    LUT4 mux_670_i25_3_lut (.A(p[24]), .B(a[24]), .C(state[0]), .Z(n1461[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i25_3_lut.init = 16'hcaca;
    LUT4 mux_670_i24_3_lut (.A(p[23]), .B(a[23]), .C(state[0]), .Z(n1461[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i24_3_lut.init = 16'hcaca;
    LUT4 mux_680_i7_3_lut (.A(csr_read_data_x[6]), .B(adder_result_x[6]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[6] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i7_3_lut.init = 16'hcaca;
    LUT4 mux_680_i8_3_lut (.A(csr_read_data_x[7]), .B(adder_result_x[7]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[7] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i8_3_lut.init = 16'hcaca;
    LUT4 mux_680_i16_3_lut (.A(csr_read_data_x[15]), .B(adder_result_x[15]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[15] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i16_3_lut.init = 16'hcaca;
    LUT4 i37703_3_lut (.A(n1562[16]), .B(n1595[16]), .C(n18869), .Z(n1793[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37703_3_lut.init = 16'hcaca;
    FD1P3AX a_i0_i15 (.D(n18918[15]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[15])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i15.GSR = "ENABLED";
    FD1P3AX cycles_19669__i5 (.D(n37[5]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(cycles[5])) /* synthesis syn_use_carry_chain=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(250[26:39])
    defparam cycles_19669__i5.GSR = "ENABLED";
    LUT4 mux_17581_i8_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[7]), 
         .C(a[6]), .D(n41417), .Z(n18884[7])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i8_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 mux_670_i23_3_lut (.A(p[22]), .B(a[22]), .C(state[0]), .Z(n1461[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i23_3_lut.init = 16'hcaca;
    LUT4 mux_670_i22_3_lut (.A(p[21]), .B(a[21]), .C(state[0]), .Z(n1461[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i22_3_lut.init = 16'hcaca;
    LUT4 i37705_3_lut (.A(n1562[15]), .B(n1595[15]), .C(n18869), .Z(n1793[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37705_3_lut.init = 16'hcaca;
    FD1P3AX a_i0_i14 (.D(n18918[14]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[14])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i14.GSR = "ENABLED";
    LUT4 mux_17581_i7_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[6]), 
         .C(a[5]), .D(n41417), .Z(n18884[6])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i7_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 mux_17581_i6_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[5]), 
         .C(a[4]), .D(n41417), .Z(n18884[5])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i6_3_lut_4_lut_4_lut.init = 16'hf0d8;
    PFUMX i27 (.BLUT(n16), .ALUT(n24948), .C0(raw_x_1), .Z(n13));
    LUT4 mux_680_i17_3_lut (.A(csr_read_data_x[16]), .B(adder_result_x[16]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[16] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i17_3_lut.init = 16'hcaca;
    LUT4 mux_680_i18_3_lut (.A(csr_read_data_x[17]), .B(adder_result_x[17]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[17] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i18_3_lut.init = 16'hcaca;
    FD1P3AX a_i0_i13 (.D(n18918[13]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[13])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i13.GSR = "ENABLED";
    FD1P3AX a_i0_i12 (.D(n18918[12]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[12])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i12.GSR = "ENABLED";
    LUT4 i21317_4_lut (.A(cycles_5__N_2497), .B(n41373), .C(divide_by_zero_x_N_2651), 
         .D(w_clk_cpu_enable_958), .Z(n23934)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i21317_4_lut.init = 16'hce0a;
    LUT4 divide_by_zero_x_I_107_4_lut (.A(cycles[3]), .B(n41408), .C(n10), 
         .D(cycles[4]), .Z(divide_by_zero_x_N_2651)) /* synthesis lut_function=(A (B)+!A (B+!(C+(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(244[17:69])
    defparam divide_by_zero_x_I_107_4_lut.init = 16'hcccd;
    LUT4 i4_4_lut (.A(cycles[2]), .B(cycles[5]), .C(cycles[0]), .D(cycles[1]), 
         .Z(n10)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(244[17:48])
    defparam i4_4_lut.init = 16'hfffe;
    LUT4 mux_17581_i5_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[4]), 
         .C(a[3]), .D(n41417), .Z(n18884[4])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i5_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 mux_680_i19_3_lut (.A(csr_read_data_x[18]), .B(adder_result_x[18]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[18] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i19_3_lut.init = 16'hcaca;
    LUT4 mux_680_i20_3_lut (.A(csr_read_data_x[19]), .B(adder_result_x[19]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[19] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i20_3_lut.init = 16'hcaca;
    LUT4 mux_17581_i4_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[3]), 
         .C(a[2]), .D(n41417), .Z(n18884[3])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i4_3_lut_4_lut_4_lut.init = 16'hf0d8;
    LUT4 mux_670_i21_3_lut (.A(p[20]), .B(a[20]), .C(state[0]), .Z(n1461[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i21_3_lut.init = 16'hcaca;
    LUT4 mux_670_i20_3_lut (.A(p[19]), .B(a[19]), .C(state[0]), .Z(n1461[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i20_3_lut.init = 16'hcaca;
    FD1P3IX b__i23 (.D(n1976[23]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[23])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i23.GSR = "ENABLED";
    LUT4 mux_17581_i3_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(bypass_data_0[2]), 
         .C(a[1]), .D(n41417), .Z(n18884[2])) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C)) */ ;
    defparam mux_17581_i3_3_lut_4_lut_4_lut.init = 16'hf0d8;
    FD1P3AX a_i0_i11 (.D(n18918[11]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[11])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i11.GSR = "ENABLED";
    LUT4 mux_680_i21_3_lut (.A(csr_read_data_x[20]), .B(adder_result_x[20]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[20] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i21_3_lut.init = 16'hcaca;
    LUT4 mux_680_i22_3_lut (.A(csr_read_data_x[21]), .B(adder_result_x[21]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[21] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i22_3_lut.init = 16'hcaca;
    LUT4 mux_680_i23_3_lut (.A(csr_read_data_x[22]), .B(adder_result_x[22]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[22] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i23_3_lut.init = 16'hcaca;
    LUT4 i29842_3_lut (.A(x_result_sel_csr_x), .B(x_result_sel_add_x), .C(x_result_sel_sext_x), 
         .Z(n24948)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i29842_3_lut.init = 16'h0101;
    LUT4 i1_4_lut (.A(n41411), .B(m_result_sel_compare_m), .C(m_result_sel_shift_m), 
         .D(direction_m), .Z(n16)) /* synthesis lut_function=(A (B+(C (D)))) */ ;
    defparam i1_4_lut.init = 16'ha888;
    LUT4 mux_697_i15_4_lut (.A(n1862[14]), .B(\instruction_d[14] ), .C(n18877), 
         .D(n41407), .Z(n1936[14])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_697_i15_4_lut.init = 16'hca0a;
    FD1P3AX a_i0_i10 (.D(n18918[10]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[10])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i10.GSR = "ENABLED";
    FD1P3IX b__i22 (.D(n1976[22]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[22])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i22.GSR = "ENABLED";
    LUT4 mux_697_i14_4_lut (.A(n1862[13]), .B(\instruction_d[13] ), .C(n18877), 
         .D(n41407), .Z(n1936[13])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_697_i14_4_lut.init = 16'hca0a;
    LUT4 mux_17583_i32_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[31]), 
         .C(n18884[31]), .D(n41417), .Z(n18918[31])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i32_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 mux_670_i19_3_lut (.A(p[18]), .B(a[18]), .C(state[0]), .Z(n1461[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i19_3_lut.init = 16'hcaca;
    LUT4 mux_670_i18_3_lut (.A(p[17]), .B(a[17]), .C(state[0]), .Z(n1461[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i18_3_lut.init = 16'hcaca;
    LUT4 mux_680_i24_3_lut (.A(csr_read_data_x[23]), .B(adder_result_x[23]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[23] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i24_3_lut.init = 16'hcaca;
    LUT4 mux_680_i25_3_lut (.A(csr_read_data_x[24]), .B(adder_result_x[24]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[24] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i25_3_lut.init = 16'hcaca;
    FD1P3IX b__i8 (.D(n1976[8]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[8])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i8.GSR = "ENABLED";
    LUT4 mux_680_i26_3_lut (.A(csr_read_data_x[25]), .B(adder_result_x[25]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[25] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i26_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_4_lut (.A(cycles_5__N_2495), .B(n42740), .C(n41364), 
         .D(n41361), .Z(n18877)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0800;
    LUT4 mux_697_i13_4_lut (.A(n1862[12]), .B(\instruction_d[12] ), .C(n18877), 
         .D(n41407), .Z(n1936[12])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_697_i13_4_lut.init = 16'hca0a;
    FD1P3AX a_i0_i9 (.D(n18918[9]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[9])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i9.GSR = "ENABLED";
    LUT4 mux_17583_i31_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[30]), 
         .C(n18884[30]), .D(n41417), .Z(n18918[30])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i31_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 mux_670_i17_3_lut (.A(p[16]), .B(a[16]), .C(state[0]), .Z(n1461[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i17_3_lut.init = 16'hcaca;
    LUT4 mux_670_i16_3_lut (.A(p[15]), .B(a[15]), .C(state[0]), .Z(n1461[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i16_3_lut.init = 16'hcaca;
    LUT4 mux_680_i27_3_lut (.A(csr_read_data_x[26]), .B(adder_result_x[26]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[26] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i27_3_lut.init = 16'hcaca;
    LUT4 mux_680_i28_3_lut (.A(csr_read_data_x[27]), .B(adder_result_x[27]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[27] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i28_3_lut.init = 16'hcaca;
    FD1P3AX a_i0_i8 (.D(n18918[8]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[8])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i8.GSR = "ENABLED";
    LUT4 mux_680_i29_3_lut (.A(csr_read_data_x[28]), .B(adder_result_x[28]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[28] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i29_3_lut.init = 16'hcaca;
    LUT4 mux_680_i1_3_lut (.A(csr_read_data_x[0]), .B(adder_result_x[0]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[0] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i1_3_lut.init = 16'hcaca;
    LUT4 mux_680_i30_3_lut (.A(csr_read_data_x[29]), .B(adder_result_x[29]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[29] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i30_3_lut.init = 16'hcaca;
    LUT4 mux_17583_i30_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[29]), 
         .C(n18884[29]), .D(n41417), .Z(n18918[29])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i30_3_lut_4_lut_4_lut.init = 16'hd8f0;
    FD1P3AX a_i0_i7 (.D(n18918[7]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[7])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i7.GSR = "ENABLED";
    LUT4 mux_17583_i29_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[28]), 
         .C(n18884[28]), .D(n41417), .Z(n18918[28])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i29_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 mux_670_i15_3_lut (.A(p[14]), .B(a[14]), .C(state[0]), .Z(n1461[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i15_3_lut.init = 16'hcaca;
    LUT4 mux_670_i14_3_lut (.A(p[13]), .B(a[13]), .C(state[0]), .Z(n1461[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i14_3_lut.init = 16'hcaca;
    FD1P3AX a_i0_i6 (.D(n18918[6]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[6])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i6.GSR = "ENABLED";
    LUT4 mux_680_i31_3_lut (.A(csr_read_data_x[30]), .B(adder_result_x[30]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[30] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i31_3_lut.init = 16'hcaca;
    LUT4 mux_680_i32_3_lut (.A(csr_read_data_x[31]), .B(adder_result_x[31]), 
         .C(x_result_sel_add_x), .Z(\x_result_31__N_616[31] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i32_3_lut.init = 16'hcaca;
    LUT4 mux_17583_i28_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[27]), 
         .C(n18884[27]), .D(n41417), .Z(n18918[27])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i28_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 mux_697_i12_4_lut (.A(n1862[11]), .B(\instruction_d[11] ), .C(n18877), 
         .D(n41407), .Z(n1936[11])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_697_i12_4_lut.init = 16'hca0a;
    LUT4 i12_3_lut_4_lut (.A(w_clk_cpu_enable_984), .B(n39970), .C(LM32I_CYC_O), 
         .D(i_cyc_o_N_1759), .Z(w_clk_cpu_enable_216)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2265[34:53])
    defparam i12_3_lut_4_lut.init = 16'hf808;
    FD1P3AX a_i0_i5 (.D(n18918[5]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[5])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i5.GSR = "ENABLED";
    FD1P3AX a_i0_i4 (.D(n18918[4]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i4.GSR = "ENABLED";
    LUT4 mux_697_i11_4_lut (.A(n1862[10]), .B(\instruction_d[10] ), .C(n18877), 
         .D(n41407), .Z(n1936[10])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_697_i11_4_lut.init = 16'hca0a;
    LUT4 mux_676_i8_3_lut (.A(operand_m[7]), .B(left_shift_result[24]), 
         .C(m_result_sel_shift_m), .Z(n1595[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i8_3_lut.init = 16'hcaca;
    LUT4 i22035_3_lut (.A(n41407), .B(\instruction_d[15] ), .C(sign_extend_immediate), 
         .Z(n24658)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i22035_3_lut.init = 16'hc4c4;
    LUT4 mux_675_i8_3_lut (.A(reg_data_1[7]), .B(w_result[7]), .C(n18863), 
         .Z(n1562[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i8_3_lut.init = 16'hcaca;
    LUT4 mux_17583_i27_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[26]), 
         .C(n18884[26]), .D(n41417), .Z(n18918[26])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i27_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 i29258_2_lut_3_lut_4_lut (.A(w_clk_cpu_enable_984), .B(n39970), 
         .C(n29[5]), .D(cycles_5__N_2495), .Z(n37[5])) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2265[34:53])
    defparam i29258_2_lut_3_lut_4_lut.init = 16'hf8f0;
    LUT4 mux_17583_i26_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[25]), 
         .C(n18884[25]), .D(n41417), .Z(n18918[25])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i26_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 mux_670_i13_3_lut (.A(p[12]), .B(a[12]), .C(state[0]), .Z(n1461[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i13_3_lut.init = 16'hcaca;
    LUT4 mux_670_i12_3_lut (.A(p[11]), .B(a[11]), .C(state[0]), .Z(n1461[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i12_3_lut.init = 16'hcaca;
    LUT4 mux_687_i32_3_lut (.A(n21414), .B(\x_result_31__N_616[31] ), .C(n18873), 
         .Z(n1862[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i32_3_lut.init = 16'hcaca;
    LUT4 mux_676_i7_3_lut (.A(operand_m[6]), .B(left_shift_result[25]), 
         .C(m_result_sel_shift_m), .Z(n1595[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i7_3_lut.init = 16'hcaca;
    LUT4 mux_675_i7_3_lut (.A(reg_data_1[6]), .B(w_result[6]), .C(n18863), 
         .Z(n1562[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i7_3_lut.init = 16'hcaca;
    FD1P3AX a_i0_i3 (.D(n18918[3]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i3.GSR = "ENABLED";
    FD1P3AX a_i0_i2 (.D(n18918[2]), .SP(w_clk_cpu_enable_865), .CK(w_clk_cpu), 
            .Q(a[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam a_i0_i2.GSR = "ENABLED";
    LUT4 mux_687_i31_3_lut (.A(n21414), .B(\x_result_31__N_616[30] ), .C(n18873), 
         .Z(n1862[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i31_3_lut.init = 16'hcaca;
    LUT4 mux_676_i6_3_lut (.A(operand_m[5]), .B(left_shift_result[26]), 
         .C(m_result_sel_shift_m), .Z(n1595[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i6_3_lut.init = 16'hcaca;
    LUT4 mux_675_i6_3_lut (.A(reg_data_1[5]), .B(w_result[5]), .C(n18863), 
         .Z(n1562[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i6_3_lut.init = 16'hcaca;
    LUT4 mux_17583_i25_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[24]), 
         .C(n18884[24]), .D(n41417), .Z(n18918[24])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i25_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 mux_17583_i24_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[23]), 
         .C(n18884[23]), .D(n41417), .Z(n18918[23])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i24_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 mux_676_i5_3_lut (.A(operand_m[4]), .B(left_shift_result[27]), 
         .C(m_result_sel_shift_m), .Z(n1595[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i5_3_lut.init = 16'hcaca;
    LUT4 mux_17583_i23_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[22]), 
         .C(n18884[22]), .D(n41417), .Z(n18918[22])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i23_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 i11_3_lut_4_lut (.A(w_clk_cpu_enable_984), .B(n39970), .C(LM32I_CYC_O), 
         .D(i_cyc_o_N_1759), .Z(n37179)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((D)+!C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2265[34:53])
    defparam i11_3_lut_4_lut.init = 16'h08f8;
    LUT4 mux_670_i11_3_lut (.A(p[10]), .B(a[10]), .C(state[0]), .Z(n1461[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i11_3_lut.init = 16'hcaca;
    LUT4 mux_670_i10_3_lut (.A(p[9]), .B(a[9]), .C(state[0]), .Z(n1461[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i10_3_lut.init = 16'hcaca;
    LUT4 mux_675_i5_3_lut (.A(reg_data_1[4]), .B(w_result[4]), .C(n18863), 
         .Z(n1562[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i5_3_lut.init = 16'hcaca;
    LUT4 mux_17583_i22_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[21]), 
         .C(n18884[21]), .D(n41417), .Z(n18918[21])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i22_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 mux_17583_i21_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[20]), 
         .C(n18884[20]), .D(n41417), .Z(n18918[20])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i21_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 mux_17583_i20_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[19]), 
         .C(n18884[19]), .D(n41417), .Z(n18918[19])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i20_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 mux_687_i30_3_lut (.A(n21414), .B(\x_result_31__N_616[29] ), .C(n18873), 
         .Z(n1862[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i30_3_lut.init = 16'hcaca;
    LUT4 mux_687_i1_3_lut (.A(\muliplicand[0] ), .B(\x_result_31__N_616[0] ), 
         .C(n18873), .Z(n1862[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i1_3_lut.init = 16'hcaca;
    LUT4 mux_670_i9_3_lut (.A(p[8]), .B(a[8]), .C(state[0]), .Z(n1461[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i9_3_lut.init = 16'hcaca;
    LUT4 mux_676_i4_3_lut (.A(operand_m[3]), .B(left_shift_result[28]), 
         .C(m_result_sel_shift_m), .Z(n1595[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i4_3_lut.init = 16'hcaca;
    LUT4 mux_670_i8_3_lut (.A(p[7]), .B(a[7]), .C(state[0]), .Z(n1461[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i8_3_lut.init = 16'hcaca;
    LUT4 mux_687_i29_3_lut (.A(n21414), .B(\x_result_31__N_616[28] ), .C(n18873), 
         .Z(n1862[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i29_3_lut.init = 16'hcaca;
    LUT4 mux_675_i4_3_lut (.A(reg_data_1[3]), .B(w_result[3]), .C(n18863), 
         .Z(n1562[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i4_3_lut.init = 16'hcaca;
    LUT4 mux_687_i28_3_lut (.A(n21414), .B(\x_result_31__N_616[27] ), .C(n18873), 
         .Z(n1862[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i28_3_lut.init = 16'hcaca;
    LUT4 mux_687_i27_3_lut (.A(n21414), .B(\x_result_31__N_616[26] ), .C(n18873), 
         .Z(n1862[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i27_3_lut.init = 16'hcaca;
    LUT4 mux_670_i1_3_lut (.A(p[0]), .B(a[0]), .C(state[0]), .Z(n1461[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i1_3_lut.init = 16'hcaca;
    LUT4 mux_17583_i19_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[18]), 
         .C(n18884[18]), .D(n41417), .Z(n18918[18])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i19_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 mux_17583_i18_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[17]), 
         .C(n18884[17]), .D(n41417), .Z(n18918[17])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i18_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 i2_4_lut_adj_273 (.A(n39272), .B(n4_adj_3775), .C(n39274), .D(n39270), 
         .Z(divide_by_zero_x_N_2647)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i2_4_lut_adj_273.init = 16'h0004;
    LUT4 i36719_4_lut (.A(b[24]), .B(n39244), .C(n39128), .D(b[30]), 
         .Z(n39272)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i36719_4_lut.init = 16'hfffe;
    LUT4 i36721_4_lut (.A(n39108), .B(n39266), .C(n39236), .D(n39104), 
         .Z(n39274)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i36721_4_lut.init = 16'hfffe;
    LUT4 mux_670_i7_3_lut (.A(p[6]), .B(a[6]), .C(state[0]), .Z(n1461[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i7_3_lut.init = 16'hcaca;
    LUT4 mux_670_i6_3_lut (.A(p[5]), .B(a[5]), .C(state[0]), .Z(n1461[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i6_3_lut.init = 16'hcaca;
    LUT4 i36717_4_lut (.A(b[1]), .B(n39240), .C(n39118), .D(b[31]), 
         .Z(n39270)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i36717_4_lut.init = 16'hfffe;
    LUT4 i36692_4_lut (.A(b[3]), .B(b[28]), .C(b[27]), .D(b[18]), .Z(n39244)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i36692_4_lut.init = 16'hfffe;
    LUT4 mux_676_i3_3_lut (.A(operand_m[2]), .B(left_shift_result[29]), 
         .C(m_result_sel_shift_m), .Z(n1595[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i3_3_lut.init = 16'hcaca;
    LUT4 mux_675_i3_3_lut (.A(reg_data_1[2]), .B(w_result[2]), .C(n18863), 
         .Z(n1562[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i3_3_lut.init = 16'hcaca;
    LUT4 mux_17583_i17_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[16]), 
         .C(n18884[16]), .D(n41417), .Z(n18918[16])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i17_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 i36581_2_lut (.A(b[2]), .B(b[5]), .Z(n39128)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i36581_2_lut.init = 16'heeee;
    LUT4 mux_687_i26_3_lut (.A(n21414), .B(\x_result_31__N_616[25] ), .C(n18873), 
         .Z(n1862[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i26_3_lut.init = 16'hcaca;
    LUT4 i36561_2_lut (.A(b[26]), .B(b[17]), .Z(n39108)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i36561_2_lut.init = 16'heeee;
    LUT4 i36713_4_lut (.A(b[22]), .B(n39232), .C(n39094), .D(b[9]), 
         .Z(n39266)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i36713_4_lut.init = 16'hfffe;
    LUT4 i36684_4_lut (.A(b[29]), .B(b[14]), .C(b[10]), .D(b[19]), .Z(n39236)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i36684_4_lut.init = 16'hfffe;
    LUT4 i36557_2_lut (.A(b[11]), .B(b[0]), .Z(n39104)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i36557_2_lut.init = 16'heeee;
    LUT4 mux_676_i2_3_lut (.A(operand_m[1]), .B(left_shift_result[30]), 
         .C(m_result_sel_shift_m), .Z(n1595[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i2_3_lut.init = 16'hcaca;
    LUT4 i36680_4_lut (.A(b[16]), .B(b[6]), .C(b[13]), .D(b[4]), .Z(n39232)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i36680_4_lut.init = 16'hfffe;
    LUT4 i36547_2_lut (.A(b[7]), .B(b[8]), .Z(n39094)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i36547_2_lut.init = 16'heeee;
    LUT4 i36688_4_lut (.A(b[20]), .B(b[21]), .C(b[12]), .D(b[25]), .Z(n39240)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i36688_4_lut.init = 16'hfffe;
    LUT4 i36571_2_lut (.A(b[23]), .B(b[15]), .Z(n39118)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i36571_2_lut.init = 16'heeee;
    LUT4 i1_3_lut (.A(cycles_5__N_2497), .B(divide_by_zero_x_N_2651), .C(state[0]), 
         .Z(n4_adj_3775)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i1_3_lut.init = 16'hc8c8;
    LUT4 mux_687_i25_3_lut (.A(n21414), .B(\x_result_31__N_616[24] ), .C(n18873), 
         .Z(n1862[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i25_3_lut.init = 16'hcaca;
    LUT4 mux_675_i2_3_lut (.A(reg_data_1[1]), .B(w_result[1]), .C(n18863), 
         .Z(n1562[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i2_3_lut.init = 16'hcaca;
    LUT4 mux_687_i24_3_lut (.A(n21414), .B(\x_result_31__N_616[23] ), .C(n18873), 
         .Z(n1862[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i24_3_lut.init = 16'hcaca;
    LUT4 mux_676_i1_3_lut (.A(operand_m[0]), .B(left_shift_result[31]), 
         .C(m_result_sel_shift_m), .Z(n1595[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i1_3_lut.init = 16'hcaca;
    LUT4 mux_670_i5_3_lut (.A(p[4]), .B(a[4]), .C(state[0]), .Z(n1461[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i5_3_lut.init = 16'hcaca;
    LUT4 mux_675_i1_3_lut (.A(reg_data_1[0]), .B(w_result[0]), .C(n18863), 
         .Z(n1562[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i1_3_lut.init = 16'hcaca;
    LUT4 mux_17583_i16_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[15]), 
         .C(n18884[15]), .D(n41417), .Z(n18918[15])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i16_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 mux_687_i23_3_lut (.A(n21414), .B(\x_result_31__N_616[22] ), .C(n18873), 
         .Z(n1862[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i23_3_lut.init = 16'hcaca;
    LUT4 mux_687_i22_3_lut (.A(n21414), .B(\x_result_31__N_616[21] ), .C(n18873), 
         .Z(n1862[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i22_3_lut.init = 16'hcaca;
    LUT4 mux_687_i21_3_lut (.A(n21414), .B(\x_result_31__N_616[20] ), .C(n18873), 
         .Z(n1862[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i21_3_lut.init = 16'hcaca;
    LUT4 mux_683_i1_3_lut (.A(n1628[0]), .B(n1285), .C(raw_x_1), .Z(n1826_c[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_683_i1_3_lut.init = 16'hcaca;
    LUT4 mux_687_i20_3_lut (.A(n21414), .B(\x_result_31__N_616[19] ), .C(n18873), 
         .Z(n1862[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i20_3_lut.init = 16'hcaca;
    LUT4 mux_687_i19_3_lut (.A(n21414), .B(\x_result_31__N_616[18] ), .C(n18873), 
         .Z(n1862[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i19_3_lut.init = 16'hcaca;
    LUT4 mux_687_i18_3_lut (.A(n21414), .B(\x_result_31__N_616[17] ), .C(n18873), 
         .Z(n1862[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i18_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_4_lut (.A(w_clk_cpu_enable_984), .B(n39970), .C(n41417), 
         .D(cycles_5__N_2495), .Z(n4)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2265[34:53])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0800;
    LUT4 mux_17583_i15_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[14]), 
         .C(n18884[14]), .D(n41417), .Z(n18918[14])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i15_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 mux_17583_i14_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[13]), 
         .C(n18884[13]), .D(n41417), .Z(n18918[13])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i14_3_lut_4_lut_4_lut.init = 16'hd8f0;
    FD1P3IX b__i21 (.D(n1976[21]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[21])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i21.GSR = "ENABLED";
    LUT4 mux_687_i17_3_lut (.A(n21414), .B(\x_result_31__N_616[16] ), .C(n18873), 
         .Z(n1862[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i17_3_lut.init = 16'hcaca;
    LUT4 mux_676_i32_3_lut (.A(operand_m[31]), .B(left_shift_result[0]), 
         .C(m_result_sel_shift_m), .Z(n1595[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i32_3_lut.init = 16'hcaca;
    LUT4 mux_675_i32_3_lut (.A(reg_data_1[31]), .B(w_result[31]), .C(n18863), 
         .Z(n1562[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i32_3_lut.init = 16'hcaca;
    LUT4 mux_676_i31_3_lut (.A(operand_m[30]), .B(left_shift_result[1]), 
         .C(m_result_sel_shift_m), .Z(n1595[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i31_3_lut.init = 16'hcaca;
    LUT4 mux_17583_i13_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[12]), 
         .C(n18884[12]), .D(n41417), .Z(n18918[12])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i13_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 mux_687_i16_3_lut (.A(n21414), .B(\x_result_31__N_616[15] ), .C(n18873), 
         .Z(n1862[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i16_3_lut.init = 16'hcaca;
    LUT4 mux_17583_i12_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[11]), 
         .C(n18884[11]), .D(n41417), .Z(n18918[11])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i12_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 mux_675_i31_3_lut (.A(reg_data_1[30]), .B(w_result[30]), .C(n18863), 
         .Z(n1562[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i31_3_lut.init = 16'hcaca;
    LUT4 mux_676_i30_3_lut (.A(operand_m[29]), .B(left_shift_result[2]), 
         .C(m_result_sel_shift_m), .Z(n1595[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i30_3_lut.init = 16'hcaca;
    LUT4 mux_687_i8_3_lut (.A(\muliplicand[7] ), .B(\x_result_31__N_616[7] ), 
         .C(n18873), .Z(n1862[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i8_3_lut.init = 16'hcaca;
    LUT4 mux_675_i30_3_lut (.A(reg_data_1[29]), .B(w_result[29]), .C(n18863), 
         .Z(n1562[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i30_3_lut.init = 16'hcaca;
    LUT4 mux_687_i7_3_lut (.A(\muliplicand[6] ), .B(\x_result_31__N_616[6] ), 
         .C(n18873), .Z(n1862[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i7_3_lut.init = 16'hcaca;
    LUT4 mux_17583_i11_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[10]), 
         .C(n18884[10]), .D(n41417), .Z(n18918[10])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i11_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 mux_676_i29_3_lut (.A(operand_m[28]), .B(left_shift_result[3]), 
         .C(m_result_sel_shift_m), .Z(n1595[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i29_3_lut.init = 16'hcaca;
    LUT4 mux_675_i29_3_lut (.A(reg_data_1[28]), .B(w_result[28]), .C(n18863), 
         .Z(n1562[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i29_3_lut.init = 16'hcaca;
    LUT4 mux_17583_i10_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[9]), 
         .C(n18884[9]), .D(n41417), .Z(n18918[9])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i10_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 mux_687_i6_3_lut (.A(\muliplicand[5] ), .B(\x_result_31__N_616[5] ), 
         .C(n18873), .Z(n1862[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i6_3_lut.init = 16'hcaca;
    LUT4 mux_676_i28_3_lut (.A(operand_m[27]), .B(left_shift_result[4]), 
         .C(m_result_sel_shift_m), .Z(n1595[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i28_3_lut.init = 16'hcaca;
    LUT4 mux_675_i28_3_lut (.A(reg_data_1[27]), .B(w_result[27]), .C(n18863), 
         .Z(n1562[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i28_3_lut.init = 16'hcaca;
    LUT4 mux_687_i5_3_lut (.A(\muliplicand[4] ), .B(\x_result_31__N_616[4] ), 
         .C(n18873), .Z(n1862[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i5_3_lut.init = 16'hcaca;
    LUT4 mux_676_i27_3_lut (.A(operand_m[26]), .B(left_shift_result[5]), 
         .C(m_result_sel_shift_m), .Z(n1595[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i27_3_lut.init = 16'hcaca;
    LUT4 mux_687_i4_3_lut (.A(\muliplicand[3] ), .B(\x_result_31__N_616[3] ), 
         .C(n18873), .Z(n1862[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i4_3_lut.init = 16'hcaca;
    FD1P3IX b__i7 (.D(n1976[7]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[7])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i7.GSR = "ENABLED";
    LUT4 i2_3_lut_4_lut_3_lut_4_lut (.A(w_clk_cpu_enable_984), .B(n39970), 
         .C(n41417), .D(cycles_5__N_2495), .Z(n22517)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2265[34:53])
    defparam i2_3_lut_4_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), 
         .C(x_result_sel_sext_x), .Z(n9)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    LUT4 i2_3_lut_4_lut_adj_274 (.A(x_result_sel_add_x), .B(x_result_sel_csr_x), 
         .C(raw_x_1), .D(n41345), .Z(n18873)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i2_3_lut_4_lut_adj_274.init = 16'he000;
    LUT4 mux_687_i3_3_lut (.A(\muliplicand[2] ), .B(\x_result_31__N_616[2] ), 
         .C(n18873), .Z(n1862[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i3_3_lut.init = 16'hcaca;
    LUT4 mux_687_i2_3_lut (.A(\muliplicand[1] ), .B(\x_result_31__N_616[1] ), 
         .C(n18873), .Z(n1862[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_687_i2_3_lut.init = 16'hcaca;
    LUT4 mux_675_i27_3_lut (.A(reg_data_1[26]), .B(w_result[26]), .C(n18863), 
         .Z(n1562[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i27_3_lut.init = 16'hcaca;
    LUT4 mux_670_i4_3_lut (.A(p[3]), .B(a[3]), .C(state[0]), .Z(n1461[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i4_3_lut.init = 16'hcaca;
    LUT4 mux_676_i26_3_lut (.A(operand_m[25]), .B(left_shift_result[6]), 
         .C(m_result_sel_shift_m), .Z(n1595[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i26_3_lut.init = 16'hcaca;
    LUT4 mux_675_i26_3_lut (.A(reg_data_1[25]), .B(w_result[25]), .C(n18863), 
         .Z(n1562[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i26_3_lut.init = 16'hcaca;
    LUT4 mux_17583_i9_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[8]), 
         .C(n18884[8]), .D(n41417), .Z(n18918[8])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i9_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 mux_676_i25_3_lut (.A(operand_m[24]), .B(left_shift_result[7]), 
         .C(m_result_sel_shift_m), .Z(n1595[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i25_3_lut.init = 16'hcaca;
    LUT4 mux_675_i25_3_lut (.A(reg_data_1[24]), .B(w_result[24]), .C(n18863), 
         .Z(n1562[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i25_3_lut.init = 16'hcaca;
    LUT4 mux_676_i24_3_lut (.A(operand_m[23]), .B(left_shift_result[8]), 
         .C(m_result_sel_shift_m), .Z(n1595[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i24_3_lut.init = 16'hcaca;
    LUT4 mux_675_i24_3_lut (.A(reg_data_1[23]), .B(w_result[23]), .C(n18863), 
         .Z(n1562[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i24_3_lut.init = 16'hcaca;
    FD1P3IX p__i31 (.D(n19597[31]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[31])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i31.GSR = "ENABLED";
    LUT4 mux_670_i3_3_lut (.A(p[2]), .B(a[2]), .C(state[0]), .Z(n1461[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_670_i3_3_lut.init = 16'hcaca;
    FD1P3IX p__i30 (.D(n19597[30]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[30])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i30.GSR = "ENABLED";
    LUT4 mux_17583_i8_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[7]), 
         .C(n18884[7]), .D(n41417), .Z(n18918[7])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i8_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 i37759_3_lut (.A(n41318), .B(n1844), .C(n18875), .Z(n1900[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37759_3_lut.init = 16'hcaca;
    LUT4 mux_676_i23_3_lut (.A(operand_m[22]), .B(left_shift_result[9]), 
         .C(m_result_sel_shift_m), .Z(n1595[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i23_3_lut.init = 16'hcaca;
    LUT4 mux_17583_i7_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[6]), 
         .C(n18884[6]), .D(n41417), .Z(n18918[6])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i7_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 mux_675_i23_3_lut (.A(reg_data_1[22]), .B(w_result[22]), .C(n18863), 
         .Z(n1562[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i23_3_lut.init = 16'hcaca;
    LUT4 mux_676_i22_3_lut (.A(operand_m[21]), .B(left_shift_result[10]), 
         .C(m_result_sel_shift_m), .Z(n1595[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i22_3_lut.init = 16'hcaca;
    LUT4 i37761_3_lut (.A(n41315), .B(n1845), .C(n18875), .Z(n1900[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37761_3_lut.init = 16'hcaca;
    LUT4 mux_675_i22_3_lut (.A(reg_data_1[21]), .B(w_result[21]), .C(n18863), 
         .Z(n1562[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i22_3_lut.init = 16'hcaca;
    FD1P3IX p__i29 (.D(n19597[29]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[29])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i29.GSR = "ENABLED";
    LUT4 mux_676_i21_3_lut (.A(operand_m[20]), .B(left_shift_result[11]), 
         .C(m_result_sel_shift_m), .Z(n1595[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i21_3_lut.init = 16'hcaca;
    LUT4 mux_675_i21_3_lut (.A(reg_data_1[20]), .B(w_result[20]), .C(n18863), 
         .Z(n1562[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i21_3_lut.init = 16'hcaca;
    LUT4 mux_676_i20_3_lut (.A(operand_m[19]), .B(left_shift_result[12]), 
         .C(m_result_sel_shift_m), .Z(n1595[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i20_3_lut.init = 16'hcaca;
    LUT4 mux_675_i20_3_lut (.A(reg_data_1[19]), .B(w_result[19]), .C(n18863), 
         .Z(n1562[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i20_3_lut.init = 16'hcaca;
    LUT4 i37763_3_lut (.A(n41307), .B(n1846), .C(n18875), .Z(n1900[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37763_3_lut.init = 16'hcaca;
    LUT4 mux_676_i19_3_lut (.A(operand_m[18]), .B(left_shift_result[13]), 
         .C(m_result_sel_shift_m), .Z(n1595[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i19_3_lut.init = 16'hcaca;
    FD1P3IX p__i28 (.D(n19597[28]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[28])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i28.GSR = "ENABLED";
    FD1P3IX p__i27 (.D(n19597[27]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[27])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i27.GSR = "ENABLED";
    LUT4 reg_data_1_10__bdd_3_lut_39268 (.A(reg_data_1[10]), .B(w_result[10]), 
         .C(n18863), .Z(n41300)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam reg_data_1_10__bdd_3_lut_39268.init = 16'hcaca;
    LUT4 reg_data_1_10__bdd_3_lut_38529 (.A(operand_m[10]), .B(m_result_sel_shift_m), 
         .C(left_shift_result[21]), .Z(n41299)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam reg_data_1_10__bdd_3_lut_38529.init = 16'he2e2;
    LUT4 i37765_3_lut (.A(n41304), .B(n1847), .C(n18875), .Z(n1900[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37765_3_lut.init = 16'hcaca;
    FD1P3IX p__i26 (.D(n19597[26]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[26])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i26.GSR = "ENABLED";
    LUT4 reg_data_1_11__bdd_3_lut_38532 (.A(operand_m[11]), .B(m_result_sel_shift_m), 
         .C(left_shift_result[20]), .Z(n41302)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam reg_data_1_11__bdd_3_lut_38532.init = 16'he2e2;
    FD1P3IX p__i25 (.D(n19597[25]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[25])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i25.GSR = "ENABLED";
    CCU2D cycles_19669_add_4_7 (.A0(cycles[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n36661), .S0(n29[5]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(250[26:39])
    defparam cycles_19669_add_4_7.INIT0 = 16'h0555;
    defparam cycles_19669_add_4_7.INIT1 = 16'h0000;
    defparam cycles_19669_add_4_7.INJECT1_0 = "NO";
    defparam cycles_19669_add_4_7.INJECT1_1 = "NO";
    LUT4 mux_675_i19_3_lut (.A(reg_data_1[18]), .B(w_result[18]), .C(n18863), 
         .Z(n1562[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_675_i19_3_lut.init = 16'hcaca;
    LUT4 mux_676_i18_3_lut (.A(operand_m[17]), .B(left_shift_result[14]), 
         .C(m_result_sel_shift_m), .Z(n1595[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_676_i18_3_lut.init = 16'hcaca;
    LUT4 reg_data_1_11__bdd_3_lut_39273 (.A(reg_data_1[11]), .B(w_result[11]), 
         .C(n18863), .Z(n41303)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam reg_data_1_11__bdd_3_lut_39273.init = 16'hcaca;
    CCU2D cycles_19669_add_4_5 (.A0(cycles[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cycles[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n36660), .COUT(n36661), .S0(n29[3]), .S1(n29[4]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(250[26:39])
    defparam cycles_19669_add_4_5.INIT0 = 16'h0555;
    defparam cycles_19669_add_4_5.INIT1 = 16'h0555;
    defparam cycles_19669_add_4_5.INJECT1_0 = "NO";
    defparam cycles_19669_add_4_5.INJECT1_1 = "NO";
    FD1P3IX p__i24 (.D(n19597[24]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[24])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i24.GSR = "ENABLED";
    FD1P3IX p__i23 (.D(n19597[23]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[23])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i23.GSR = "ENABLED";
    LUT4 reg_data_1_12__bdd_3_lut_38535 (.A(operand_m[12]), .B(m_result_sel_shift_m), 
         .C(left_shift_result[19]), .Z(n41305)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam reg_data_1_12__bdd_3_lut_38535.init = 16'he2e2;
    CCU2D cycles_19669_add_4_3 (.A0(cycles[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cycles[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n36659), .COUT(n36660), .S0(n29[1]), .S1(n29[2]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(250[26:39])
    defparam cycles_19669_add_4_3.INIT0 = 16'h0555;
    defparam cycles_19669_add_4_3.INIT1 = 16'h0555;
    defparam cycles_19669_add_4_3.INJECT1_0 = "NO";
    defparam cycles_19669_add_4_3.INJECT1_1 = "NO";
    LUT4 reg_data_1_12__bdd_3_lut_39278 (.A(reg_data_1[12]), .B(w_result[12]), 
         .C(n18863), .Z(n41306)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam reg_data_1_12__bdd_3_lut_39278.init = 16'hcaca;
    LUT4 i37687_3_lut (.A(n1562[24]), .B(n1595[24]), .C(n18869), .Z(n1793[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37687_3_lut.init = 16'hcaca;
    FD1P3IX p__i22 (.D(n19597[22]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[22])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i22.GSR = "ENABLED";
    FD1P3IX p__i21 (.D(n19597[21]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[21])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i21.GSR = "ENABLED";
    LUT4 mux_697_i10_4_lut (.A(n1862[9]), .B(\instruction_d[9] ), .C(n18877), 
         .D(n41407), .Z(n1936[9])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_697_i10_4_lut.init = 16'hca0a;
    FD1P3IX p__i20 (.D(n19597[20]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[20])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i20.GSR = "ENABLED";
    FD1P3IX p__i19 (.D(n19597[19]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[19])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i19.GSR = "ENABLED";
    CCU2D cycles_19669_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cycles[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n36659), .S1(n29[0]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(250[26:39])
    defparam cycles_19669_add_4_1.INIT0 = 16'hF000;
    defparam cycles_19669_add_4_1.INIT1 = 16'h0555;
    defparam cycles_19669_add_4_1.INJECT1_0 = "NO";
    defparam cycles_19669_add_4_1.INJECT1_1 = "NO";
    LUT4 mux_697_i9_4_lut (.A(n1862[8]), .B(\instruction_d[8] ), .C(n18877), 
         .D(n41407), .Z(n1936[8])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_697_i9_4_lut.init = 16'hca0a;
    FD1P3IX p__i18 (.D(n19597[18]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[18])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i18.GSR = "ENABLED";
    FD1P3IX p__i17 (.D(n19597[17]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[17])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i17.GSR = "ENABLED";
    LUT4 reg_data_1_13__bdd_3_lut_38541 (.A(operand_m[13]), .B(m_result_sel_shift_m), 
         .C(left_shift_result[18]), .Z(n41313)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam reg_data_1_13__bdd_3_lut_38541.init = 16'he2e2;
    LUT4 reg_data_1_13__bdd_3_lut_39283 (.A(reg_data_1[13]), .B(w_result[13]), 
         .C(n18863), .Z(n41314)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam reg_data_1_13__bdd_3_lut_39283.init = 16'hcaca;
    LUT4 i37650_3_lut (.A(n1562[7]), .B(n1595[7]), .C(n18869), .Z(n1793[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37650_3_lut.init = 16'hcaca;
    LUT4 i21323_4_lut (.A(cycles_5__N_2495), .B(n4_adj_3775), .C(n42740), 
         .D(n38799), .Z(n23940)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i21323_4_lut.init = 16'heece;
    FD1P3IX p__i16 (.D(n19597[16]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[16])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i16.GSR = "ENABLED";
    LUT4 reg_data_1_14__bdd_3_lut_38544 (.A(operand_m[14]), .B(m_result_sel_shift_m), 
         .C(left_shift_result[17]), .Z(n41316)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam reg_data_1_14__bdd_3_lut_38544.init = 16'he2e2;
    FD1P3IX p__i15 (.D(n19597[15]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[15])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i15.GSR = "ENABLED";
    LUT4 reg_data_1_14__bdd_3_lut_39289 (.A(reg_data_1[14]), .B(w_result[14]), 
         .C(n18863), .Z(n41317)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam reg_data_1_14__bdd_3_lut_39289.init = 16'hcaca;
    PFUMX i38128 (.BLUT(n40483), .ALUT(n40482), .C0(n18869), .Z(n40484));
    LUT4 i21321_3_lut (.A(state[0]), .B(n38840), .C(divide_by_zero_x_N_2651), 
         .Z(n23938)) /* synthesis lut_function=(A (B+!(C))+!A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i21321_3_lut.init = 16'hcece;
    FD1P3IX p__i14 (.D(n19597[14]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[14])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i14.GSR = "ENABLED";
    LUT4 i37652_3_lut (.A(n1562[6]), .B(n1595[6]), .C(n18869), .Z(n1793[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37652_3_lut.init = 16'hcaca;
    LUT4 mux_17583_i6_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[5]), 
         .C(n18884[5]), .D(n41417), .Z(n18918[5])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i6_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 mux_17583_i5_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[4]), 
         .C(n18884[4]), .D(n41417), .Z(n18918[4])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i5_3_lut_4_lut_4_lut.init = 16'hd8f0;
    FD1P3IX p__i13 (.D(n19597[13]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[13])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i13.GSR = "ENABLED";
    LUT4 i37654_3_lut (.A(n1562[5]), .B(n1595[5]), .C(n18869), .Z(n1793[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37654_3_lut.init = 16'hcaca;
    FD1P3IX p__i12 (.D(n19597[12]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[12])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i12.GSR = "ENABLED";
    FD1P3IX p__i11 (.D(n19597[11]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[11])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i11.GSR = "ENABLED";
    L6MUX21 mux_705_i2 (.D0(n1900[1]), .D1(n1936[1]), .SD(n18879), .Z(n1976[1]));
    L6MUX21 mux_705_i3 (.D0(n1900[2]), .D1(n1936[2]), .SD(n18879), .Z(n1976[2]));
    PFUMX i38123 (.BLUT(n40477), .ALUT(n40476), .C0(n18869), .Z(n40478));
    FD1P3IX p__i10 (.D(n19597[10]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[10])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i10.GSR = "ENABLED";
    L6MUX21 mux_705_i4 (.D0(n1900[3]), .D1(n1936[3]), .SD(n18879), .Z(n1976[3]));
    FD1P3IX p__i9 (.D(n19597[9]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[9])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i9.GSR = "ENABLED";
    LUT4 i37656_3_lut (.A(n1562[4]), .B(n1595[4]), .C(n18869), .Z(n1793[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37656_3_lut.init = 16'hcaca;
    L6MUX21 mux_705_i5 (.D0(n1900[4]), .D1(n1936[4]), .SD(n18879), .Z(n1976[4]));
    L6MUX21 mux_705_i6 (.D0(n1900[5]), .D1(n1936[5]), .SD(n18879), .Z(n1976[5]));
    L6MUX21 mux_705_i7 (.D0(n1900[6]), .D1(n1936[6]), .SD(n18879), .Z(n1976[6]));
    L6MUX21 mux_705_i8 (.D0(n1900[7]), .D1(n1936[7]), .SD(n18879), .Z(n1976[7]));
    PFUMX mux_705_i9 (.BLUT(n1900[8]), .ALUT(n1936[8]), .C0(n18879), .Z(n1976[8]));
    LUT4 i37658_3_lut (.A(n1562[3]), .B(n1595[3]), .C(n18869), .Z(n1793[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37658_3_lut.init = 16'hcaca;
    PFUMX mux_705_i10 (.BLUT(n1900[9]), .ALUT(n1936[9]), .C0(n18879), 
          .Z(n1976[9]));
    FD1P3IX p__i8 (.D(n19597[8]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[8])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i8.GSR = "ENABLED";
    LUT4 i37660_3_lut (.A(n1562[2]), .B(n1595[2]), .C(n18869), .Z(n1793[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37660_3_lut.init = 16'hcaca;
    FD1P3IX p__i7 (.D(n19597[7]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[7])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i7.GSR = "ENABLED";
    PFUMX mux_705_i11 (.BLUT(n1900[10]), .ALUT(n1936[10]), .C0(n18879), 
          .Z(n1976[10]));
    LUT4 i37662_3_lut (.A(n1562[1]), .B(n1595[1]), .C(n18869), .Z(n1793[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37662_3_lut.init = 16'hcaca;
    L6MUX21 mux_705_i1 (.D0(n1900[0]), .D1(n1936[0]), .SD(n18879), .Z(n1976[0]));
    PFUMX mux_705_i12 (.BLUT(n1900[11]), .ALUT(n1936[11]), .C0(n18879), 
          .Z(n1976[11]));
    PFUMX mux_705_i13 (.BLUT(n1900[12]), .ALUT(n1936[12]), .C0(n18879), 
          .Z(n1976[12]));
    FD1P3AX result_x_i0_i31 (.D(n1461[31]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[31])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i31.GSR = "ENABLED";
    FD1P3IX p__i6 (.D(n19597[6]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[6])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i6.GSR = "ENABLED";
    FD1P3IX p__i5 (.D(n19597[5]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[5])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i5.GSR = "ENABLED";
    PFUMX mux_705_i14 (.BLUT(n1900[13]), .ALUT(n1936[13]), .C0(n18879), 
          .Z(n1976[13]));
    LUT4 mux_17583_i4_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[3]), 
         .C(n18884[3]), .D(n41417), .Z(n18918[3])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i4_3_lut_4_lut_4_lut.init = 16'hd8f0;
    LUT4 mux_17583_i3_3_lut_4_lut_4_lut (.A(w_clk_cpu_enable_958), .B(pc_f[2]), 
         .C(n18884[2]), .D(n41417), .Z(n18918[2])) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A (C)) */ ;
    defparam mux_17583_i3_3_lut_4_lut_4_lut.init = 16'hd8f0;
    PFUMX mux_705_i15 (.BLUT(n1900[14]), .ALUT(n1936[14]), .C0(n18879), 
          .Z(n1976[14]));
    LUT4 i37664_3_lut (.A(n1562[0]), .B(n1595[0]), .C(n18869), .Z(n1793[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37664_3_lut.init = 16'hcaca;
    LUT4 mux_680_i15_3_lut (.A(csr_read_data_x[14]), .B(adder_result_x[14]), 
         .C(x_result_sel_add_x), .Z(n1727[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i15_3_lut.init = 16'hcaca;
    L6MUX21 mux_705_i16 (.D0(n1900[15]), .D1(n1936[15]), .SD(n18879), 
            .Z(n1976[15]));
    L6MUX21 mux_705_i17 (.D0(n1900[16]), .D1(n1936[16]), .SD(n18879), 
            .Z(n1976[16]));
    FD1P3AX result_x_i0_i30 (.D(n1461[30]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[30])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i30.GSR = "ENABLED";
    FD1P3AX result_x_i0_i29 (.D(n1461[29]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[29])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i29.GSR = "ENABLED";
    FD1P3IX p__i4 (.D(n19597[4]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i4.GSR = "ENABLED";
    LUT4 mux_680_i14_3_lut (.A(csr_read_data_x[13]), .B(adder_result_x[13]), 
         .C(x_result_sel_add_x), .Z(n1727[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i14_3_lut.init = 16'hcaca;
    FD1P3IX p__i3 (.D(n19597[3]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i3.GSR = "ENABLED";
    L6MUX21 mux_705_i18 (.D0(n1900[17]), .D1(n1936[17]), .SD(n18879), 
            .Z(n1976[17]));
    L6MUX21 mux_705_i19 (.D0(n1900[18]), .D1(n1936[18]), .SD(n18879), 
            .Z(n1976[18]));
    L6MUX21 mux_705_i20 (.D0(n1900[19]), .D1(n1936[19]), .SD(n18879), 
            .Z(n1976[19]));
    L6MUX21 mux_705_i21 (.D0(n1900[20]), .D1(n1936[20]), .SD(n18879), 
            .Z(n1976[20]));
    LUT4 mux_680_i13_3_lut (.A(csr_read_data_x[12]), .B(adder_result_x[12]), 
         .C(x_result_sel_add_x), .Z(n1727[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i13_3_lut.init = 16'hcaca;
    L6MUX21 mux_705_i22 (.D0(n1900[21]), .D1(n1936[21]), .SD(n18879), 
            .Z(n1976[21]));
    L6MUX21 mux_705_i23 (.D0(n1900[22]), .D1(n1936[22]), .SD(n18879), 
            .Z(n1976[22]));
    L6MUX21 mux_705_i24 (.D0(n1900[23]), .D1(n1936[23]), .SD(n18879), 
            .Z(n1976[23]));
    L6MUX21 mux_705_i25 (.D0(n1900[24]), .D1(n1936[24]), .SD(n18879), 
            .Z(n1976[24]));
    L6MUX21 mux_705_i26 (.D0(n1900[25]), .D1(n1936[25]), .SD(n18879), 
            .Z(n1976[25]));
    L6MUX21 mux_705_i27 (.D0(n1900[26]), .D1(n1936[26]), .SD(n18879), 
            .Z(n1976[26]));
    L6MUX21 mux_705_i28 (.D0(n1900[27]), .D1(n1936[27]), .SD(n18879), 
            .Z(n1976[27]));
    L6MUX21 mux_705_i29 (.D0(n1900[28]), .D1(n1936[28]), .SD(n18879), 
            .Z(n1976[28]));
    L6MUX21 mux_705_i30 (.D0(n1900[29]), .D1(n1936[29]), .SD(n18879), 
            .Z(n1976[29]));
    L6MUX21 mux_705_i31 (.D0(n1900[30]), .D1(n1936[30]), .SD(n18879), 
            .Z(n1976[30]));
    L6MUX21 mux_705_i32 (.D0(n1900[31]), .D1(n1936[31]), .SD(n18879), 
            .Z(n1976[31]));
    FD1P3AX result_x_i0_i28 (.D(n1461[28]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[28])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i28.GSR = "ENABLED";
    FD1P3AX result_x_i0_i27 (.D(n1461[27]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[27])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i27.GSR = "ENABLED";
    FD1P3IX p__i2 (.D(n19597[2]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i2.GSR = "ENABLED";
    FD1P3IX p__i1 (.D(n19597[1]), .SP(w_clk_cpu_enable_865), .CD(w_clk_cpu_enable_958), 
            .CK(w_clk_cpu), .Q(p[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam p__i1.GSR = "ENABLED";
    PFUMX mux_697_i2 (.BLUT(n1862[1]), .ALUT(n1791), .C0(n18877), .Z(n1936[1]));
    CCU2D p_30__I_0_add_2_33 (.A0(p[30]), .B0(b[31]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n36651), 
          .S0(t[31]), .S1(t[32]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam p_30__I_0_add_2_33.INIT0 = 16'h5999;
    defparam p_30__I_0_add_2_33.INIT1 = 16'hffff;
    defparam p_30__I_0_add_2_33.INJECT1_0 = "NO";
    defparam p_30__I_0_add_2_33.INJECT1_1 = "NO";
    PFUMX mux_697_i3 (.BLUT(n1862[2]), .ALUT(n1790), .C0(n18877), .Z(n1936[2]));
    FD1P3AX result_x_i0_i26 (.D(n1461[26]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[26])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i26.GSR = "ENABLED";
    FD1P3AX result_x_i0_i25 (.D(n1461[25]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[25])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i25.GSR = "ENABLED";
    PFUMX mux_697_i4 (.BLUT(n1862[3]), .ALUT(n1789), .C0(n18877), .Z(n1936[3]));
    LUT4 mux_680_i12_3_lut (.A(csr_read_data_x[11]), .B(adder_result_x[11]), 
         .C(x_result_sel_add_x), .Z(n1727[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i12_3_lut.init = 16'hcaca;
    LUT4 mux_680_i11_3_lut (.A(csr_read_data_x[10]), .B(adder_result_x[10]), 
         .C(x_result_sel_add_x), .Z(n1727[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i11_3_lut.init = 16'hcaca;
    PFUMX mux_697_i5 (.BLUT(n1862[4]), .ALUT(n1788), .C0(n18877), .Z(n1936[4]));
    PFUMX mux_697_i6 (.BLUT(n1862[5]), .ALUT(n1787), .C0(n18877), .Z(n1936[5]));
    LUT4 mux_680_i10_3_lut (.A(csr_read_data_x[9]), .B(adder_result_x[9]), 
         .C(x_result_sel_add_x), .Z(n1727[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i10_3_lut.init = 16'hcaca;
    FD1P3AX result_x_i0_i24 (.D(n1461[24]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[24])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i24.GSR = "ENABLED";
    FD1P3AX result_x_i0_i23 (.D(n1461[23]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[23])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i23.GSR = "ENABLED";
    PFUMX mux_697_i7 (.BLUT(n1862[6]), .ALUT(n1786), .C0(n18877), .Z(n1936[6]));
    PFUMX mux_697_i8 (.BLUT(n1862[7]), .ALUT(n1785), .C0(n18877), .Z(n1936[7]));
    LUT4 mux_680_i9_3_lut (.A(csr_read_data_x[8]), .B(adder_result_x[8]), 
         .C(x_result_sel_add_x), .Z(n1727[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam mux_680_i9_3_lut.init = 16'hcaca;
    PFUMX mux_697_i16 (.BLUT(n1862[15]), .ALUT(n1777), .C0(n18877), .Z(n1936[15]));
    LUT4 i37673_3_lut (.A(n1562[31]), .B(n1595[31]), .C(n18869), .Z(n1793[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37673_3_lut.init = 16'hcaca;
    LUT4 i37675_3_lut (.A(n1562[30]), .B(n1595[30]), .C(n18869), .Z(n1793[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37675_3_lut.init = 16'hcaca;
    CCU2D p_30__I_0_add_2_31 (.A0(p[28]), .B0(b[29]), .C0(GND_net), .D0(GND_net), 
          .A1(p[29]), .B1(b[30]), .C1(GND_net), .D1(GND_net), .CIN(n36650), 
          .COUT(n36651), .S0(t[29]), .S1(t[30]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam p_30__I_0_add_2_31.INIT0 = 16'h5999;
    defparam p_30__I_0_add_2_31.INIT1 = 16'h5999;
    defparam p_30__I_0_add_2_31.INJECT1_0 = "NO";
    defparam p_30__I_0_add_2_31.INJECT1_1 = "NO";
    FD1P3AX result_x_i0_i22 (.D(n1461[22]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[22])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i22.GSR = "ENABLED";
    FD1P3AX result_x_i0_i21 (.D(n1461[21]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[21])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i21.GSR = "ENABLED";
    LUT4 i37685_3_lut (.A(n1562[25]), .B(n1595[25]), .C(n18869), .Z(n1793[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37685_3_lut.init = 16'hcaca;
    PFUMX mux_697_i17 (.BLUT(n1862[16]), .ALUT(n1776), .C0(n18877), .Z(n1936[16]));
    CCU2D p_30__I_0_add_2_29 (.A0(p[26]), .B0(b[27]), .C0(GND_net), .D0(GND_net), 
          .A1(p[27]), .B1(b[28]), .C1(GND_net), .D1(GND_net), .CIN(n36649), 
          .COUT(n36650), .S0(t[27]), .S1(t[28]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam p_30__I_0_add_2_29.INIT0 = 16'h5999;
    defparam p_30__I_0_add_2_29.INIT1 = 16'h5999;
    defparam p_30__I_0_add_2_29.INJECT1_0 = "NO";
    defparam p_30__I_0_add_2_29.INJECT1_1 = "NO";
    CCU2D p_30__I_0_add_2_27 (.A0(p[24]), .B0(b[25]), .C0(GND_net), .D0(GND_net), 
          .A1(p[25]), .B1(b[26]), .C1(GND_net), .D1(GND_net), .CIN(n36648), 
          .COUT(n36649), .S0(t[25]), .S1(t[26]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam p_30__I_0_add_2_27.INIT0 = 16'h5999;
    defparam p_30__I_0_add_2_27.INIT1 = 16'h5999;
    defparam p_30__I_0_add_2_27.INJECT1_0 = "NO";
    defparam p_30__I_0_add_2_27.INJECT1_1 = "NO";
    PFUMX mux_697_i18 (.BLUT(n1862[17]), .ALUT(n1775), .C0(n18877), .Z(n1936[17]));
    LUT4 i37677_3_lut (.A(n1562[29]), .B(n1595[29]), .C(n18869), .Z(n1793[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37677_3_lut.init = 16'hcaca;
    PFUMX mux_697_i19 (.BLUT(n1862[18]), .ALUT(n1774), .C0(n18877), .Z(n1936[18]));
    PFUMX mux_697_i20 (.BLUT(n1862[19]), .ALUT(n1773), .C0(n18877), .Z(n1936[19]));
    FD1P3AX result_x_i0_i20 (.D(n1461[20]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[20])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i20.GSR = "ENABLED";
    FD1P3AX result_x_i0_i19 (.D(n1461[19]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[19])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i19.GSR = "ENABLED";
    CCU2D p_30__I_0_add_2_25 (.A0(p[22]), .B0(b[23]), .C0(GND_net), .D0(GND_net), 
          .A1(p[23]), .B1(b[24]), .C1(GND_net), .D1(GND_net), .CIN(n36647), 
          .COUT(n36648), .S0(t[23]), .S1(t[24]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam p_30__I_0_add_2_25.INIT0 = 16'h5999;
    defparam p_30__I_0_add_2_25.INIT1 = 16'h5999;
    defparam p_30__I_0_add_2_25.INJECT1_0 = "NO";
    defparam p_30__I_0_add_2_25.INJECT1_1 = "NO";
    CCU2D p_30__I_0_add_2_23 (.A0(p[20]), .B0(b[21]), .C0(GND_net), .D0(GND_net), 
          .A1(p[21]), .B1(b[22]), .C1(GND_net), .D1(GND_net), .CIN(n36646), 
          .COUT(n36647), .S0(t[21]), .S1(t[22]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam p_30__I_0_add_2_23.INIT0 = 16'h5999;
    defparam p_30__I_0_add_2_23.INIT1 = 16'h5999;
    defparam p_30__I_0_add_2_23.INJECT1_0 = "NO";
    defparam p_30__I_0_add_2_23.INJECT1_1 = "NO";
    LUT4 i37679_3_lut (.A(n1562[28]), .B(n1595[28]), .C(n18869), .Z(n1793[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37679_3_lut.init = 16'hcaca;
    PFUMX mux_697_i21 (.BLUT(n1862[20]), .ALUT(n1772), .C0(n18877), .Z(n1936[20]));
    PFUMX mux_697_i22 (.BLUT(n1862[21]), .ALUT(n1771), .C0(n18877), .Z(n1936[21]));
    PFUMX mux_697_i23 (.BLUT(n1862[22]), .ALUT(n1770), .C0(n18877), .Z(n1936[22]));
    FD1P3AX result_x_i0_i18 (.D(n1461[18]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[18])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i18.GSR = "ENABLED";
    LUT4 i37681_3_lut (.A(n1562[27]), .B(n1595[27]), .C(n18869), .Z(n1793[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37681_3_lut.init = 16'hcaca;
    FD1P3AX result_x_i0_i17 (.D(n1461[17]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[17])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i17.GSR = "ENABLED";
    PFUMX mux_697_i24 (.BLUT(n1862[23]), .ALUT(n1769), .C0(n18877), .Z(n1936[23]));
    PFUMX mux_697_i25 (.BLUT(n1862[24]), .ALUT(n1768), .C0(n18877), .Z(n1936[24]));
    PFUMX mux_697_i26 (.BLUT(n1862[25]), .ALUT(n1767), .C0(n18877), .Z(n1936[25]));
    FD1P3AX result_x_i0_i16 (.D(n1461[16]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[16])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i16.GSR = "ENABLED";
    FD1P3AX result_x_i0_i15 (.D(n1461[15]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[15])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i15.GSR = "ENABLED";
    CCU2D p_30__I_0_add_2_21 (.A0(p[18]), .B0(b[19]), .C0(GND_net), .D0(GND_net), 
          .A1(p[19]), .B1(b[20]), .C1(GND_net), .D1(GND_net), .CIN(n36645), 
          .COUT(n36646), .S0(t[19]), .S1(t[20]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam p_30__I_0_add_2_21.INIT0 = 16'h5999;
    defparam p_30__I_0_add_2_21.INIT1 = 16'h5999;
    defparam p_30__I_0_add_2_21.INJECT1_0 = "NO";
    defparam p_30__I_0_add_2_21.INJECT1_1 = "NO";
    CCU2D p_30__I_0_add_2_19 (.A0(p[16]), .B0(b[17]), .C0(GND_net), .D0(GND_net), 
          .A1(p[17]), .B1(b[18]), .C1(GND_net), .D1(GND_net), .CIN(n36644), 
          .COUT(n36645), .S0(t[17]), .S1(t[18]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam p_30__I_0_add_2_19.INIT0 = 16'h5999;
    defparam p_30__I_0_add_2_19.INIT1 = 16'h5999;
    defparam p_30__I_0_add_2_19.INJECT1_0 = "NO";
    defparam p_30__I_0_add_2_19.INJECT1_1 = "NO";
    CCU2D p_30__I_0_add_2_17 (.A0(p[14]), .B0(b[15]), .C0(GND_net), .D0(GND_net), 
          .A1(p[15]), .B1(b[16]), .C1(GND_net), .D1(GND_net), .CIN(n36643), 
          .COUT(n36644), .S0(t[15]), .S1(t[16]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam p_30__I_0_add_2_17.INIT0 = 16'h5999;
    defparam p_30__I_0_add_2_17.INIT1 = 16'h5999;
    defparam p_30__I_0_add_2_17.INJECT1_0 = "NO";
    defparam p_30__I_0_add_2_17.INJECT1_1 = "NO";
    PFUMX mux_697_i27 (.BLUT(n1862[26]), .ALUT(n1766), .C0(n18877), .Z(n1936[26]));
    PFUMX mux_697_i28 (.BLUT(n1862[27]), .ALUT(n1765), .C0(n18877), .Z(n1936[27]));
    PFUMX mux_697_i29 (.BLUT(n1862[28]), .ALUT(n1764), .C0(n18877), .Z(n1936[28]));
    PFUMX mux_697_i1 (.BLUT(n1862[0]), .ALUT(n1792), .C0(n18877), .Z(n1936[0]));
    PFUMX mux_697_i30 (.BLUT(n1862[29]), .ALUT(n1763), .C0(n18877), .Z(n1936[29]));
    FD1P3AX result_x_i0_i14 (.D(n1461[14]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[14])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i14.GSR = "ENABLED";
    FD1P3AX result_x_i0_i13 (.D(n1461[13]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[13])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i13.GSR = "ENABLED";
    CCU2D p_30__I_0_add_2_15 (.A0(p[12]), .B0(b[13]), .C0(GND_net), .D0(GND_net), 
          .A1(p[13]), .B1(b[14]), .C1(GND_net), .D1(GND_net), .CIN(n36642), 
          .COUT(n36643), .S0(t[13]), .S1(t[14]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam p_30__I_0_add_2_15.INIT0 = 16'h5999;
    defparam p_30__I_0_add_2_15.INIT1 = 16'h5999;
    defparam p_30__I_0_add_2_15.INJECT1_0 = "NO";
    defparam p_30__I_0_add_2_15.INJECT1_1 = "NO";
    PFUMX mux_697_i31 (.BLUT(n1862[30]), .ALUT(n1762), .C0(n18877), .Z(n1936[30]));
    PFUMX mux_697_i32 (.BLUT(n1862[31]), .ALUT(n24658), .C0(n18877), .Z(n1936[31]));
    FD1P3AX result_x_i0_i12 (.D(n1461[12]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[12])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i12.GSR = "ENABLED";
    FD1P3AX result_x_i0_i11 (.D(n1461[11]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[11])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i11.GSR = "ENABLED";
    CCU2D p_30__I_0_add_2_13 (.A0(p[10]), .B0(b[11]), .C0(GND_net), .D0(GND_net), 
          .A1(p[11]), .B1(b[12]), .C1(GND_net), .D1(GND_net), .CIN(n36641), 
          .COUT(n36642), .S0(t[11]), .S1(t[12]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam p_30__I_0_add_2_13.INIT0 = 16'h5999;
    defparam p_30__I_0_add_2_13.INIT1 = 16'h5999;
    defparam p_30__I_0_add_2_13.INJECT1_0 = "NO";
    defparam p_30__I_0_add_2_13.INJECT1_1 = "NO";
    CCU2D p_30__I_0_add_2_11 (.A0(p[8]), .B0(b[9]), .C0(GND_net), .D0(GND_net), 
          .A1(p[9]), .B1(b[10]), .C1(GND_net), .D1(GND_net), .CIN(n36640), 
          .COUT(n36641), .S0(t[9]), .S1(t[10]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam p_30__I_0_add_2_11.INIT0 = 16'h5999;
    defparam p_30__I_0_add_2_11.INIT1 = 16'h5999;
    defparam p_30__I_0_add_2_11.INJECT1_0 = "NO";
    defparam p_30__I_0_add_2_11.INJECT1_1 = "NO";
    CCU2D p_30__I_0_add_2_9 (.A0(p[6]), .B0(b[7]), .C0(GND_net), .D0(GND_net), 
          .A1(p[7]), .B1(b[8]), .C1(GND_net), .D1(GND_net), .CIN(n36639), 
          .COUT(n36640), .S0(t[7]), .S1(t[8]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(156[12:64])
    defparam p_30__I_0_add_2_9.INIT0 = 16'h5999;
    defparam p_30__I_0_add_2_9.INIT1 = 16'h5999;
    defparam p_30__I_0_add_2_9.INJECT1_0 = "NO";
    defparam p_30__I_0_add_2_9.INJECT1_1 = "NO";
    FD1P3AX result_x_i0_i10 (.D(n1461[10]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[10])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i10.GSR = "ENABLED";
    FD1P3AX result_x_i0_i9 (.D(n1461[9]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[9])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i9.GSR = "ENABLED";
    LUT4 i37683_3_lut (.A(n1562[26]), .B(n1595[26]), .C(n18869), .Z(n1793[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(191[9] 305[16])
    defparam i37683_3_lut.init = 16'hcaca;
    PFUMX mux_693_i16 (.BLUT(n1793[15]), .ALUT(n1843), .C0(n18875), .Z(n1900[15]));
    PFUMX mux_693_i17 (.BLUT(n1793[16]), .ALUT(n1842), .C0(n18875), .Z(n1900[16]));
    FD1P3IX b__i6 (.D(n1976[6]), .SP(w_clk_cpu_enable_958), .CD(n22517), 
            .CK(w_clk_cpu), .Q(b[6])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam b__i6.GSR = "ENABLED";
    FD1P3AX result_x_i0_i8 (.D(n1461[8]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[8])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i8.GSR = "ENABLED";
    FD1P3AX result_x_i0_i7 (.D(n1461[7]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[7])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i7.GSR = "ENABLED";
    PFUMX mux_693_i18 (.BLUT(n1793[17]), .ALUT(n1841), .C0(n18875), .Z(n1900[17]));
    PFUMX mux_693_i19 (.BLUT(n1793[18]), .ALUT(n1840), .C0(n18875), .Z(n1900[18]));
    PFUMX mux_693_i20 (.BLUT(n1793[19]), .ALUT(n1839), .C0(n18875), .Z(n1900[19]));
    FD1P3AX result_x_i0_i6 (.D(n1461[6]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[6])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i6.GSR = "ENABLED";
    FD1P3AX result_x_i0_i5 (.D(n1461[5]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[5])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i5.GSR = "ENABLED";
    PFUMX mux_693_i21 (.BLUT(n1793[20]), .ALUT(n1838), .C0(n18875), .Z(n1900[20]));
    PFUMX mux_693_i22 (.BLUT(n1793[21]), .ALUT(n1837), .C0(n18875), .Z(n1900[21]));
    FD1P3AX result_x_i0_i4 (.D(n1461[4]), .SP(mc_stall_request_x), .CK(w_clk_cpu), 
            .Q(mc_result_x[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=20, LSE_RCOL=6, LSE_LLINE=1102, LSE_RLINE=1128 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_mc_arithmetic.v(187[5] 306[8])
    defparam result_x_i0_i4.GSR = "ENABLED";
    PFUMX mux_693_i23 (.BLUT(n1793[22]), .ALUT(n1836), .C0(n18875), .Z(n1900[22]));
    PFUMX mux_693_i24 (.BLUT(n1793[23]), .ALUT(n1835), .C0(n18875), .Z(n1900[23]));
    
endmodule
//
// Verilog Description of module lm32_logic_op
//

module lm32_logic_op (\logic_op_x[2] , \logic_op_x[3] , muliplicand, \condition_x[0] , 
            \size_x[1] , operand_1_x, logic_result_x) /* synthesis syn_module_defined=1 */ ;
    input \logic_op_x[2] ;
    input \logic_op_x[3] ;
    input [31:0]muliplicand;
    input \condition_x[0] ;
    input \size_x[1] ;
    input [31:0]operand_1_x;
    output [31:0]logic_result_x;
    
    
    wire n39713, n39712, n39710, n39709, n39707, n39706, n39704, 
        n39703, n39701, n39700, n39698, n39697, n39695, n39694, 
        n39692, n39691, n39689, n39688, n39686, n39685, n39683, 
        n39682, n39680, n39679, n39677, n39676, n39674, n39673, 
        n39671, n39670, n39668, n39667, n39665, n39664, n39662, 
        n39661, n39659, n39658, n39656, n39655, n39749, n39748, 
        n39746, n39745, n39743, n39742, n39740, n39739, n39737, 
        n39736, n39734, n39733, n39731, n39730, n39728, n39727, 
        n39725, n39724, n39722, n39721, n39719, n39718, n39716, 
        n39715;
    
    LUT4 i37159_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[13]), 
         .Z(n39713)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37159_3_lut.init = 16'hcaca;
    LUT4 i37158_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[13]), 
         .Z(n39712)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37158_3_lut.init = 16'hcaca;
    LUT4 i37156_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[14]), 
         .Z(n39710)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37156_3_lut.init = 16'hcaca;
    LUT4 i37155_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[14]), 
         .Z(n39709)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37155_3_lut.init = 16'hcaca;
    LUT4 i37153_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[15]), 
         .Z(n39707)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37153_3_lut.init = 16'hcaca;
    LUT4 i37152_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[15]), 
         .Z(n39706)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37152_3_lut.init = 16'hcaca;
    LUT4 i37150_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[16]), 
         .Z(n39704)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37150_3_lut.init = 16'hcaca;
    LUT4 i37149_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[16]), 
         .Z(n39703)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37149_3_lut.init = 16'hcaca;
    LUT4 i37147_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[17]), 
         .Z(n39701)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37147_3_lut.init = 16'hcaca;
    LUT4 i37146_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[17]), 
         .Z(n39700)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37146_3_lut.init = 16'hcaca;
    LUT4 i37144_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[18]), 
         .Z(n39698)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37144_3_lut.init = 16'hcaca;
    LUT4 i37143_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[18]), 
         .Z(n39697)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37143_3_lut.init = 16'hcaca;
    LUT4 i37141_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[19]), 
         .Z(n39695)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37141_3_lut.init = 16'hcaca;
    LUT4 i37140_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[19]), 
         .Z(n39694)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37140_3_lut.init = 16'hcaca;
    LUT4 i37138_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[20]), 
         .Z(n39692)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37138_3_lut.init = 16'hcaca;
    LUT4 i37137_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[20]), 
         .Z(n39691)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37137_3_lut.init = 16'hcaca;
    LUT4 i37135_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[21]), 
         .Z(n39689)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37135_3_lut.init = 16'hcaca;
    LUT4 i37134_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[21]), 
         .Z(n39688)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37134_3_lut.init = 16'hcaca;
    LUT4 i37132_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[22]), 
         .Z(n39686)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37132_3_lut.init = 16'hcaca;
    LUT4 i37131_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[22]), 
         .Z(n39685)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37131_3_lut.init = 16'hcaca;
    LUT4 i37129_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[23]), 
         .Z(n39683)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37129_3_lut.init = 16'hcaca;
    LUT4 i37128_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[23]), 
         .Z(n39682)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37128_3_lut.init = 16'hcaca;
    LUT4 i37126_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[24]), 
         .Z(n39680)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37126_3_lut.init = 16'hcaca;
    LUT4 i37125_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[24]), 
         .Z(n39679)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37125_3_lut.init = 16'hcaca;
    LUT4 i37123_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[25]), 
         .Z(n39677)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37123_3_lut.init = 16'hcaca;
    LUT4 i37122_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[25]), 
         .Z(n39676)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37122_3_lut.init = 16'hcaca;
    LUT4 i37120_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[26]), 
         .Z(n39674)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37120_3_lut.init = 16'hcaca;
    LUT4 i37119_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[26]), 
         .Z(n39673)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37119_3_lut.init = 16'hcaca;
    LUT4 i37117_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[27]), 
         .Z(n39671)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37117_3_lut.init = 16'hcaca;
    LUT4 i37116_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[27]), 
         .Z(n39670)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37116_3_lut.init = 16'hcaca;
    LUT4 i37114_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[28]), 
         .Z(n39668)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37114_3_lut.init = 16'hcaca;
    LUT4 i37113_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[28]), 
         .Z(n39667)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37113_3_lut.init = 16'hcaca;
    LUT4 i37111_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[29]), 
         .Z(n39665)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37111_3_lut.init = 16'hcaca;
    LUT4 i37110_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[29]), 
         .Z(n39664)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37110_3_lut.init = 16'hcaca;
    LUT4 i37108_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[0]), 
         .Z(n39662)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37108_3_lut.init = 16'hcaca;
    LUT4 i37107_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[0]), 
         .Z(n39661)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37107_3_lut.init = 16'hcaca;
    LUT4 i37105_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[30]), 
         .Z(n39659)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37105_3_lut.init = 16'hcaca;
    LUT4 i37104_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[30]), 
         .Z(n39658)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37104_3_lut.init = 16'hcaca;
    LUT4 i37102_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[31]), 
         .Z(n39656)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37102_3_lut.init = 16'hcaca;
    LUT4 i37101_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[31]), 
         .Z(n39655)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37101_3_lut.init = 16'hcaca;
    LUT4 i37195_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[1]), 
         .Z(n39749)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37195_3_lut.init = 16'hcaca;
    LUT4 i37194_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[1]), 
         .Z(n39748)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37194_3_lut.init = 16'hcaca;
    LUT4 i37192_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[2]), 
         .Z(n39746)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37192_3_lut.init = 16'hcaca;
    LUT4 i37191_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[2]), 
         .Z(n39745)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37191_3_lut.init = 16'hcaca;
    LUT4 i37189_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[3]), 
         .Z(n39743)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37189_3_lut.init = 16'hcaca;
    LUT4 i37188_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[3]), 
         .Z(n39742)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37188_3_lut.init = 16'hcaca;
    LUT4 i37186_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[4]), 
         .Z(n39740)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37186_3_lut.init = 16'hcaca;
    LUT4 i37185_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[4]), 
         .Z(n39739)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37185_3_lut.init = 16'hcaca;
    LUT4 i37183_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[5]), 
         .Z(n39737)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37183_3_lut.init = 16'hcaca;
    LUT4 i37182_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[5]), 
         .Z(n39736)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37182_3_lut.init = 16'hcaca;
    LUT4 i37180_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[6]), 
         .Z(n39734)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37180_3_lut.init = 16'hcaca;
    LUT4 i37179_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[6]), 
         .Z(n39733)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37179_3_lut.init = 16'hcaca;
    LUT4 i37177_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[7]), 
         .Z(n39731)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37177_3_lut.init = 16'hcaca;
    LUT4 i37176_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[7]), 
         .Z(n39730)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37176_3_lut.init = 16'hcaca;
    LUT4 i37174_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[8]), 
         .Z(n39728)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37174_3_lut.init = 16'hcaca;
    LUT4 i37173_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[8]), 
         .Z(n39727)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37173_3_lut.init = 16'hcaca;
    LUT4 i37171_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[9]), 
         .Z(n39725)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37171_3_lut.init = 16'hcaca;
    LUT4 i37170_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[9]), 
         .Z(n39724)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37170_3_lut.init = 16'hcaca;
    LUT4 i37168_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[10]), 
         .Z(n39722)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37168_3_lut.init = 16'hcaca;
    LUT4 i37167_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[10]), 
         .Z(n39721)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37167_3_lut.init = 16'hcaca;
    LUT4 i37165_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[11]), 
         .Z(n39719)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37165_3_lut.init = 16'hcaca;
    LUT4 i37164_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[11]), 
         .Z(n39718)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37164_3_lut.init = 16'hcaca;
    LUT4 i37162_3_lut (.A(\logic_op_x[2] ), .B(\logic_op_x[3] ), .C(muliplicand[12]), 
         .Z(n39716)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37162_3_lut.init = 16'hcaca;
    LUT4 i37161_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(muliplicand[12]), 
         .Z(n39715)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i37161_3_lut.init = 16'hcaca;
    PFUMX i37103 (.BLUT(n39655), .ALUT(n39656), .C0(operand_1_x[31]), 
          .Z(logic_result_x[31]));
    PFUMX i37106 (.BLUT(n39658), .ALUT(n39659), .C0(operand_1_x[30]), 
          .Z(logic_result_x[30]));
    PFUMX i37109 (.BLUT(n39661), .ALUT(n39662), .C0(operand_1_x[0]), .Z(logic_result_x[0]));
    PFUMX i37112 (.BLUT(n39664), .ALUT(n39665), .C0(operand_1_x[29]), 
          .Z(logic_result_x[29]));
    PFUMX i37115 (.BLUT(n39667), .ALUT(n39668), .C0(operand_1_x[28]), 
          .Z(logic_result_x[28]));
    PFUMX i37118 (.BLUT(n39670), .ALUT(n39671), .C0(operand_1_x[27]), 
          .Z(logic_result_x[27]));
    PFUMX i37121 (.BLUT(n39673), .ALUT(n39674), .C0(operand_1_x[26]), 
          .Z(logic_result_x[26]));
    PFUMX i37124 (.BLUT(n39676), .ALUT(n39677), .C0(operand_1_x[25]), 
          .Z(logic_result_x[25]));
    PFUMX i37127 (.BLUT(n39679), .ALUT(n39680), .C0(operand_1_x[24]), 
          .Z(logic_result_x[24]));
    PFUMX i37130 (.BLUT(n39682), .ALUT(n39683), .C0(operand_1_x[23]), 
          .Z(logic_result_x[23]));
    PFUMX i37133 (.BLUT(n39685), .ALUT(n39686), .C0(operand_1_x[22]), 
          .Z(logic_result_x[22]));
    PFUMX i37136 (.BLUT(n39688), .ALUT(n39689), .C0(operand_1_x[21]), 
          .Z(logic_result_x[21]));
    PFUMX i37139 (.BLUT(n39691), .ALUT(n39692), .C0(operand_1_x[20]), 
          .Z(logic_result_x[20]));
    PFUMX i37142 (.BLUT(n39694), .ALUT(n39695), .C0(operand_1_x[19]), 
          .Z(logic_result_x[19]));
    PFUMX i37145 (.BLUT(n39697), .ALUT(n39698), .C0(operand_1_x[18]), 
          .Z(logic_result_x[18]));
    PFUMX i37148 (.BLUT(n39700), .ALUT(n39701), .C0(operand_1_x[17]), 
          .Z(logic_result_x[17]));
    PFUMX i37151 (.BLUT(n39703), .ALUT(n39704), .C0(operand_1_x[16]), 
          .Z(logic_result_x[16]));
    PFUMX i37154 (.BLUT(n39706), .ALUT(n39707), .C0(operand_1_x[15]), 
          .Z(logic_result_x[15]));
    PFUMX i37157 (.BLUT(n39709), .ALUT(n39710), .C0(operand_1_x[14]), 
          .Z(logic_result_x[14]));
    PFUMX i37160 (.BLUT(n39712), .ALUT(n39713), .C0(operand_1_x[13]), 
          .Z(logic_result_x[13]));
    PFUMX i37163 (.BLUT(n39715), .ALUT(n39716), .C0(operand_1_x[12]), 
          .Z(logic_result_x[12]));
    PFUMX i37166 (.BLUT(n39718), .ALUT(n39719), .C0(operand_1_x[11]), 
          .Z(logic_result_x[11]));
    PFUMX i37169 (.BLUT(n39721), .ALUT(n39722), .C0(operand_1_x[10]), 
          .Z(logic_result_x[10]));
    PFUMX i37172 (.BLUT(n39724), .ALUT(n39725), .C0(operand_1_x[9]), .Z(logic_result_x[9]));
    PFUMX i37175 (.BLUT(n39727), .ALUT(n39728), .C0(operand_1_x[8]), .Z(logic_result_x[8]));
    PFUMX i37178 (.BLUT(n39730), .ALUT(n39731), .C0(operand_1_x[7]), .Z(logic_result_x[7]));
    PFUMX i37181 (.BLUT(n39733), .ALUT(n39734), .C0(operand_1_x[6]), .Z(logic_result_x[6]));
    PFUMX i37184 (.BLUT(n39736), .ALUT(n39737), .C0(operand_1_x[5]), .Z(logic_result_x[5]));
    PFUMX i37187 (.BLUT(n39739), .ALUT(n39740), .C0(operand_1_x[4]), .Z(logic_result_x[4]));
    PFUMX i37190 (.BLUT(n39742), .ALUT(n39743), .C0(operand_1_x[3]), .Z(logic_result_x[3]));
    PFUMX i37193 (.BLUT(n39745), .ALUT(n39746), .C0(operand_1_x[2]), .Z(logic_result_x[2]));
    PFUMX i37196 (.BLUT(n39748), .ALUT(n39749), .C0(operand_1_x[1]), .Z(logic_result_x[1]));
    
endmodule
//
// Verilog Description of module lm32_load_store_unit
//

module lm32_load_store_unit (store_operand_x, \condition_x[0] , \size_x[1] , 
            wb_load_complete, w_clk_cpu, w_clk_cpu_enable_972, LM32D_WE_O, 
            w_clk_cpu_enable_886, n41372, LM32D_DAT_O, w_clk_cpu_enable_623, 
            SHAREDBUS_DAT_O, LM32D_ADR_O, operand_m, LM32D_SEL_O, LM32D_STB_O, 
            w_clk_cpu_enable_245, n41492, byte_enable_x, LM32D_CYC_O, 
            n26096, n26122, \operand_w[0] , load_data_w, \operand_w[1] , 
            n2, n2_adj_49, \byte_enable_x[1] , wb_load_complete_N_2129, 
            w_clk_cpu_enable_711, stall_wb_load_N_2112, n42746, n46, 
            n4, n41428, n41491, \adder_result_x[1] , \adder_result_x[0] , 
            wb_select_m, w_clk_cpu_enable_878, n42726, \store_data_x[31] , 
            \store_data_x[30] , sign_extend_x, w_clk_cpu_enable_985, \store_data_x[15] , 
            stall_wb_load, exception_m, \store_data_x[14] ) /* synthesis syn_module_defined=1 */ ;
    input [31:0]store_operand_x;
    input \condition_x[0] ;
    input \size_x[1] ;
    output wb_load_complete;
    input w_clk_cpu;
    input w_clk_cpu_enable_972;
    output LM32D_WE_O;
    input w_clk_cpu_enable_886;
    input n41372;
    output [31:0]LM32D_DAT_O;
    input w_clk_cpu_enable_623;
    input [31:0]SHAREDBUS_DAT_O;
    output [31:0]LM32D_ADR_O;
    input [31:0]operand_m;
    output [3:0]LM32D_SEL_O;
    output LM32D_STB_O;
    input w_clk_cpu_enable_245;
    input n41492;
    input [3:0]byte_enable_x;
    output LM32D_CYC_O;
    input n26096;
    input n26122;
    input \operand_w[0] ;
    output [31:0]load_data_w;
    input \operand_w[1] ;
    output n2;
    output n2_adj_49;
    input \byte_enable_x[1] ;
    input wb_load_complete_N_2129;
    input w_clk_cpu_enable_711;
    input stall_wb_load_N_2112;
    input n42746;
    input n46;
    input n4;
    input n41428;
    input n41491;
    input \adder_result_x[1] ;
    input \adder_result_x[0] ;
    output wb_select_m;
    input w_clk_cpu_enable_878;
    input n42726;
    input \store_data_x[31] ;
    input \store_data_x[30] ;
    input sign_extend_x;
    input w_clk_cpu_enable_985;
    input \store_data_x[15] ;
    output stall_wb_load;
    input exception_m;
    input \store_data_x[14] ;
    
    wire w_clk_cpu /* synthesis SET_AS_NETWORK=w_clk_cpu, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(22[6:15])
    wire [31:0]store_data_x;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(243[22:34])
    
    wire n2_c, n2_adj_3699, n2_adj_3700, w_clk_cpu_enable_27, d_we_o_N_2124;
    wire [31:0]store_data_m;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(244[22:34])
    
    wire n2_adj_3701;
    wire [1:0]size_m;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(239[22:28])
    wire [31:0]data_m;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(247[23:29])
    
    wire w_clk_cpu_enable_438;
    wire [3:0]byte_enable_m;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(246[29:42])
    wire [1:0]size_w;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(240[22:28])
    wire [31:0]data_w;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(248[22:28])
    
    wire sign_extend_w, sign_extend_m, n30, n28, n31, n41506, n41505, 
        n35, n32, n27, n32_adj_3702, n32_adj_3703, n32_adj_3704, 
        n32_adj_3705, n23, n28_adj_3706, n31_adj_3707, n32_adj_3709, 
        n25, n25_adj_3711, n36, n2_adj_3712, n25_adj_3713, n25_adj_3714, 
        n25_adj_3715, n25_adj_3716, n2_adj_3717, n25_adj_3718, n32_adj_3719, 
        n32_adj_3720;
    wire [3:0]byte_enable_x_c;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(245[29:42])
    
    wire n11, n11_adj_3721, n11_adj_3722, n11_adj_3723, n11_adj_3724, 
        n11_adj_3725, n11_adj_3726, n17, n32_adj_3727, n32_adj_3728, 
        n32_adj_3729, n32_adj_3730, n36_adj_3731, n32_adj_3732, n32_adj_3733, 
        n31_adj_3734, n31_adj_3735, n31_adj_3736, n36_adj_3737, n36_adj_3738, 
        n36_adj_3739, n36_adj_3740, n36_adj_3741, n33, n36_adj_3742, 
        n33_adj_3743, n31_adj_3744, n31_adj_3745, n31_adj_3746, w_clk_cpu_enable_979, 
        n32_adj_3747, n32_adj_3748, n23_adj_3749, n28_adj_3750, n23_adj_3751, 
        n28_adj_3752, n23_adj_3753, n28_adj_3754, n23_adj_3755, n28_adj_3756, 
        n23_adj_3757, n28_adj_3758, n23_adj_3759, n28_adj_3760, n32389;
    
    LUT4 size_x_1__I_0_153_Mux_10_i3_3_lut_4_lut (.A(store_operand_x[2]), 
         .B(\condition_x[0] ), .C(\size_x[1] ), .D(store_operand_x[10]), 
         .Z(store_data_x[10])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_153_Mux_10_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_153_Mux_26_i3_3_lut_4_lut (.A(store_operand_x[2]), 
         .B(\condition_x[0] ), .C(\size_x[1] ), .D(n2_c), .Z(store_data_x[26])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_153_Mux_26_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_153_Mux_11_i3_3_lut_4_lut (.A(store_operand_x[3]), 
         .B(\condition_x[0] ), .C(\size_x[1] ), .D(store_operand_x[11]), 
         .Z(store_data_x[11])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_153_Mux_11_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_153_Mux_27_i3_3_lut_4_lut (.A(store_operand_x[3]), 
         .B(\condition_x[0] ), .C(\size_x[1] ), .D(n2_adj_3699), .Z(store_data_x[27])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_153_Mux_27_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_153_Mux_12_i3_3_lut_4_lut (.A(store_operand_x[4]), 
         .B(\condition_x[0] ), .C(\size_x[1] ), .D(store_operand_x[12]), 
         .Z(store_data_x[12])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_153_Mux_12_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_153_Mux_28_i3_3_lut_4_lut (.A(store_operand_x[4]), 
         .B(\condition_x[0] ), .C(\size_x[1] ), .D(n2_adj_3700), .Z(store_data_x[28])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_153_Mux_28_i3_3_lut_4_lut.init = 16'hf202;
    FD1P3IX wb_load_complete_135 (.D(d_we_o_N_2124), .SP(w_clk_cpu_enable_27), 
            .CD(w_clk_cpu_enable_972), .CK(w_clk_cpu), .Q(wb_load_complete));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_load_complete_135.GSR = "ENABLED";
    FD1P3AX store_data_m_i0_i13 (.D(store_data_x[13]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(store_data_m[13])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i13.GSR = "ENABLED";
    FD1P3AX store_data_m_i0_i12 (.D(store_data_x[12]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(store_data_m[12])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i12.GSR = "ENABLED";
    FD1P3AX store_data_m_i0_i11 (.D(store_data_x[11]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(store_data_m[11])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i11.GSR = "ENABLED";
    FD1P3AX store_data_m_i0_i10 (.D(store_data_x[10]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(store_data_m[10])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i10.GSR = "ENABLED";
    LUT4 size_x_1__I_0_153_Mux_13_i3_3_lut_4_lut (.A(store_operand_x[5]), 
         .B(\condition_x[0] ), .C(\size_x[1] ), .D(store_operand_x[13]), 
         .Z(store_data_x[13])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_153_Mux_13_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_153_Mux_29_i3_3_lut_4_lut (.A(store_operand_x[5]), 
         .B(\condition_x[0] ), .C(\size_x[1] ), .D(n2_adj_3701), .Z(store_data_x[29])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_153_Mux_29_i3_3_lut_4_lut.init = 16'hf202;
    FD1P3AX store_data_m_i0_i9 (.D(store_data_x[9]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(store_data_m[9])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i9.GSR = "ENABLED";
    FD1P3AX store_data_m_i0_i8 (.D(store_data_x[8]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(store_data_m[8])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i8.GSR = "ENABLED";
    FD1P3AX size_m_i0_i0 (.D(\condition_x[0] ), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(size_m[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam size_m_i0_i0.GSR = "ENABLED";
    FD1P3AX d_we_o_130 (.D(n41372), .SP(w_clk_cpu_enable_886), .CK(w_clk_cpu), 
            .Q(LM32D_WE_O));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_we_o_130.GSR = "ENABLED";
    FD1P3AX d_dat_o_i0_i0 (.D(store_data_m[0]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i0.GSR = "ENABLED";
    FD1P3AX wb_data_m_i0_i0 (.D(SHAREDBUS_DAT_O[0]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i0.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i0 (.D(operand_m[0]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i0.GSR = "ENABLED";
    FD1P3AX d_sel_o_i0_i0 (.D(byte_enable_m[0]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_SEL_O[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_sel_o_i0_i0.GSR = "ENABLED";
    FD1P3AX d_stb_o_126 (.D(n41492), .SP(w_clk_cpu_enable_245), .CK(w_clk_cpu), 
            .Q(LM32D_STB_O)) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_stb_o_126.GSR = "ENABLED";
    FD1P3AX byte_enable_m_i0_i0 (.D(byte_enable_x[0]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(byte_enable_m[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam byte_enable_m_i0_i0.GSR = "ENABLED";
    FD1S3AX size_w_i0 (.D(size_m[0]), .CK(w_clk_cpu), .Q(size_w[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam size_w_i0.GSR = "ENABLED";
    FD1S3AX data_w_i0 (.D(data_m[0]), .CK(w_clk_cpu), .Q(data_w[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i0.GSR = "ENABLED";
    FD1S3AX sign_extend_w_144 (.D(sign_extend_m), .CK(w_clk_cpu), .Q(sign_extend_w)) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam sign_extend_w_144.GSR = "ENABLED";
    FD1S3AX d_cyc_o_125 (.D(n26096), .CK(w_clk_cpu), .Q(LM32D_CYC_O)) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_cyc_o_125.GSR = "ENABLED";
    FD1P3IX store_data_m_i0_i1 (.D(store_operand_x[1]), .SP(w_clk_cpu_enable_972), 
            .CD(n26122), .CK(w_clk_cpu), .Q(store_data_m[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i1.GSR = "ENABLED";
    PFUMX i44 (.BLUT(n30), .ALUT(n28), .C0(\operand_w[0] ), .Z(n31));
    LUT4 i1_4_lut (.A(sign_extend_w), .B(n41506), .C(n41505), .D(\operand_w[0] ), 
         .Z(n35)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(527[22:31])
    defparam i1_4_lut.init = 16'ha088;
    LUT4 i55_3_lut (.A(n32), .B(n27), .C(size_w[0]), .Z(load_data_w[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut.init = 16'hcaca;
    LUT4 i55_3_lut_adj_192 (.A(n32_adj_3702), .B(n27), .C(size_w[0]), 
         .Z(load_data_w[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_192.init = 16'hcaca;
    LUT4 i55_3_lut_adj_193 (.A(n32_adj_3703), .B(n27), .C(size_w[0]), 
         .Z(load_data_w[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_193.init = 16'hcaca;
    LUT4 i55_3_lut_adj_194 (.A(n32_adj_3704), .B(n27), .C(size_w[0]), 
         .Z(load_data_w[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_194.init = 16'hcaca;
    LUT4 i55_3_lut_adj_195 (.A(n32_adj_3705), .B(n27), .C(size_w[0]), 
         .Z(load_data_w[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_195.init = 16'hcaca;
    FD1P3AX wb_data_m_i0_i31 (.D(SHAREDBUS_DAT_O[31]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[31])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i31.GSR = "ENABLED";
    FD1P3AX wb_data_m_i0_i30 (.D(SHAREDBUS_DAT_O[30]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[30])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i30.GSR = "ENABLED";
    FD1P3AX wb_data_m_i0_i29 (.D(SHAREDBUS_DAT_O[29]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[29])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i29.GSR = "ENABLED";
    FD1P3AX wb_data_m_i0_i28 (.D(SHAREDBUS_DAT_O[28]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[28])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i28.GSR = "ENABLED";
    FD1P3AX wb_data_m_i0_i27 (.D(SHAREDBUS_DAT_O[27]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[27])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i27.GSR = "ENABLED";
    FD1P3AX wb_data_m_i0_i26 (.D(SHAREDBUS_DAT_O[26]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[26])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i26.GSR = "ENABLED";
    FD1P3AX wb_data_m_i0_i25 (.D(SHAREDBUS_DAT_O[25]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[25])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i25.GSR = "ENABLED";
    FD1P3AX wb_data_m_i0_i24 (.D(SHAREDBUS_DAT_O[24]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[24])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i24.GSR = "ENABLED";
    PFUMX i52 (.BLUT(n23), .ALUT(n28_adj_3706), .C0(\operand_w[1] ), .Z(n31_adj_3707));
    FD1P3AX wb_data_m_i0_i23 (.D(SHAREDBUS_DAT_O[23]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[23])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i23.GSR = "ENABLED";
    FD1P3AX wb_data_m_i0_i22 (.D(SHAREDBUS_DAT_O[22]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[22])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i22.GSR = "ENABLED";
    LUT4 size_x_1__I_0_153_Mux_31_i2_3_lut (.A(store_operand_x[31]), .B(store_operand_x[15]), 
         .C(\condition_x[0] ), .Z(n2)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_153_Mux_31_i2_3_lut.init = 16'hcaca;
    LUT4 i55_3_lut_adj_196 (.A(n32_adj_3709), .B(n27), .C(size_w[0]), 
         .Z(load_data_w[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_196.init = 16'hcaca;
    FD1P3AX wb_data_m_i0_i21 (.D(SHAREDBUS_DAT_O[21]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[21])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i21.GSR = "ENABLED";
    FD1P3AX wb_data_m_i0_i20 (.D(SHAREDBUS_DAT_O[20]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[20])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i20.GSR = "ENABLED";
    FD1P3AX wb_data_m_i0_i19 (.D(SHAREDBUS_DAT_O[19]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[19])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i19.GSR = "ENABLED";
    FD1P3AX wb_data_m_i0_i18 (.D(SHAREDBUS_DAT_O[18]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[18])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i18.GSR = "ENABLED";
    FD1P3AX wb_data_m_i0_i17 (.D(SHAREDBUS_DAT_O[17]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[17])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i17.GSR = "ENABLED";
    FD1P3AX wb_data_m_i0_i16 (.D(SHAREDBUS_DAT_O[16]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[16])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i16.GSR = "ENABLED";
    LUT4 size_x_1__I_0_153_Mux_30_i2_3_lut (.A(store_operand_x[30]), .B(store_operand_x[14]), 
         .C(\condition_x[0] ), .Z(n2_adj_49)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_153_Mux_30_i2_3_lut.init = 16'hcaca;
    FD1P3AX wb_data_m_i0_i15 (.D(SHAREDBUS_DAT_O[15]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[15])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i15.GSR = "ENABLED";
    FD1P3AX wb_data_m_i0_i14 (.D(SHAREDBUS_DAT_O[14]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[14])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i14.GSR = "ENABLED";
    LUT4 store_operand_x_0__bdd_4_lut (.A(store_operand_x[0]), .B(\size_x[1] ), 
         .C(store_operand_x[16]), .D(\condition_x[0] ), .Z(store_data_x[16])) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(((D)+!C)+!B)) */ ;
    defparam store_operand_x_0__bdd_4_lut.init = 16'h88e2;
    LUT4 size_x_1__I_0_153_Mux_29_i2_3_lut (.A(store_operand_x[29]), .B(store_operand_x[13]), 
         .C(\condition_x[0] ), .Z(n2_adj_3701)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_153_Mux_29_i2_3_lut.init = 16'hcaca;
    LUT4 size_x_1__I_0_153_Mux_28_i2_3_lut (.A(store_operand_x[28]), .B(store_operand_x[12]), 
         .C(\condition_x[0] ), .Z(n2_adj_3700)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_153_Mux_28_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut (.A(data_w[18]), .B(data_w[2]), .C(\operand_w[1] ), 
         .D(size_w[0]), .Z(n25)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut.init = 16'hcacc;
    FD1P3AX wb_data_m_i0_i13 (.D(SHAREDBUS_DAT_O[13]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[13])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i13.GSR = "ENABLED";
    FD1P3AX wb_data_m_i0_i12 (.D(SHAREDBUS_DAT_O[12]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[12])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i12.GSR = "ENABLED";
    LUT4 size_x_1__I_0_153_Mux_27_i2_3_lut (.A(store_operand_x[27]), .B(store_operand_x[11]), 
         .C(\condition_x[0] ), .Z(n2_adj_3699)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_153_Mux_27_i2_3_lut.init = 16'hcaca;
    FD1P3AX wb_data_m_i0_i11 (.D(SHAREDBUS_DAT_O[11]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[11])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i11.GSR = "ENABLED";
    FD1P3AX wb_data_m_i0_i10 (.D(SHAREDBUS_DAT_O[10]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[10])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i10.GSR = "ENABLED";
    LUT4 size_x_1__I_0_153_Mux_26_i2_3_lut (.A(store_operand_x[26]), .B(store_operand_x[10]), 
         .C(\condition_x[0] ), .Z(n2_c)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_153_Mux_26_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut_adj_197 (.A(data_w[17]), .B(data_w[1]), .C(\operand_w[1] ), 
         .D(size_w[0]), .Z(n25_adj_3711)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_197.init = 16'hcacc;
    LUT4 i51_4_lut_4_lut (.A(size_w[0]), .B(\operand_w[1] ), .C(data_w[7]), 
         .D(data_w[23]), .Z(n36)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam i51_4_lut_4_lut.init = 16'hf2d0;
    LUT4 store_operand_x_1__bdd_4_lut (.A(store_operand_x[1]), .B(\size_x[1] ), 
         .C(store_operand_x[17]), .D(\condition_x[0] ), .Z(store_data_x[17])) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(((D)+!C)+!B)) */ ;
    defparam store_operand_x_1__bdd_4_lut.init = 16'h88e2;
    FD1P3AX wb_data_m_i0_i9 (.D(SHAREDBUS_DAT_O[9]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[9])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i9.GSR = "ENABLED";
    FD1P3AX wb_data_m_i0_i8 (.D(SHAREDBUS_DAT_O[8]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[8])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i8.GSR = "ENABLED";
    LUT4 size_x_1__I_0_153_Mux_25_i2_3_lut (.A(store_operand_x[25]), .B(store_operand_x[9]), 
         .C(\condition_x[0] ), .Z(n2_adj_3712)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_153_Mux_25_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut_adj_198 (.A(data_w[22]), .B(data_w[6]), .C(\operand_w[1] ), 
         .D(size_w[0]), .Z(n25_adj_3713)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_198.init = 16'hcacc;
    LUT4 i1_4_lut_4_lut_adj_199 (.A(data_w[21]), .B(data_w[5]), .C(\operand_w[1] ), 
         .D(size_w[0]), .Z(n25_adj_3714)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_199.init = 16'hcacc;
    FD1P3AX wb_data_m_i0_i7 (.D(SHAREDBUS_DAT_O[7]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[7])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i7.GSR = "ENABLED";
    FD1P3AX wb_data_m_i0_i6 (.D(SHAREDBUS_DAT_O[6]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[6])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i6.GSR = "ENABLED";
    LUT4 i1_4_lut_4_lut_adj_200 (.A(data_w[20]), .B(data_w[4]), .C(\operand_w[1] ), 
         .D(size_w[0]), .Z(n25_adj_3715)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_200.init = 16'hcacc;
    LUT4 i1_4_lut_4_lut_adj_201 (.A(data_w[16]), .B(data_w[0]), .C(\operand_w[1] ), 
         .D(size_w[0]), .Z(n25_adj_3716)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_201.init = 16'hcacc;
    LUT4 size_x_1__I_0_153_Mux_24_i2_3_lut (.A(store_operand_x[24]), .B(store_operand_x[8]), 
         .C(\condition_x[0] ), .Z(n2_adj_3717)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_153_Mux_24_i2_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut_adj_202 (.A(data_w[19]), .B(data_w[3]), .C(\operand_w[1] ), 
         .D(size_w[0]), .Z(n25_adj_3718)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_202.init = 16'hcacc;
    FD1P3AX wb_data_m_i0_i5 (.D(SHAREDBUS_DAT_O[5]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[5])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i5.GSR = "ENABLED";
    FD1P3AX wb_data_m_i0_i4 (.D(SHAREDBUS_DAT_O[4]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i4.GSR = "ENABLED";
    LUT4 i55_3_lut_adj_203 (.A(n32_adj_3719), .B(n27), .C(size_w[0]), 
         .Z(load_data_w[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_203.init = 16'hcaca;
    FD1P3AX wb_data_m_i0_i3 (.D(SHAREDBUS_DAT_O[3]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i3.GSR = "ENABLED";
    FD1P3AX wb_data_m_i0_i2 (.D(SHAREDBUS_DAT_O[2]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i2.GSR = "ENABLED";
    LUT4 i55_3_lut_adj_204 (.A(n32_adj_3720), .B(n27), .C(size_w[0]), 
         .Z(load_data_w[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_204.init = 16'hcaca;
    FD1P3AX wb_data_m_i0_i1 (.D(SHAREDBUS_DAT_O[1]), .SP(w_clk_cpu_enable_438), 
            .CK(w_clk_cpu), .Q(data_m[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam wb_data_m_i0_i1.GSR = "ENABLED";
    FD1P3AX d_dat_o_i0_i31 (.D(store_data_m[31]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[31])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i31.GSR = "ENABLED";
    FD1P3AX byte_enable_m_i0_i3 (.D(byte_enable_x_c[3]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(byte_enable_m[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam byte_enable_m_i0_i3.GSR = "ENABLED";
    LUT4 i2_2_lut_3_lut (.A(\operand_w[1] ), .B(size_w[0]), .C(data_w[24]), 
         .Z(n11)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i2_2_lut_3_lut.init = 16'h4040;
    LUT4 i2_2_lut_3_lut_adj_205 (.A(\operand_w[1] ), .B(size_w[0]), .C(data_w[25]), 
         .Z(n11_adj_3721)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i2_2_lut_3_lut_adj_205.init = 16'h4040;
    LUT4 i2_2_lut_3_lut_adj_206 (.A(\operand_w[1] ), .B(size_w[0]), .C(data_w[27]), 
         .Z(n11_adj_3722)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i2_2_lut_3_lut_adj_206.init = 16'h4040;
    FD1P3AX d_dat_o_i0_i30 (.D(store_data_m[30]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[30])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i30.GSR = "ENABLED";
    FD1P3AX d_dat_o_i0_i29 (.D(store_data_m[29]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[29])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i29.GSR = "ENABLED";
    FD1P3AX byte_enable_m_i0_i2 (.D(byte_enable_x_c[2]), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(byte_enable_m[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam byte_enable_m_i0_i2.GSR = "ENABLED";
    LUT4 i2_2_lut_3_lut_adj_207 (.A(\operand_w[1] ), .B(size_w[0]), .C(data_w[26]), 
         .Z(n11_adj_3723)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i2_2_lut_3_lut_adj_207.init = 16'h4040;
    LUT4 i2_2_lut_3_lut_adj_208 (.A(\operand_w[1] ), .B(size_w[0]), .C(data_w[28]), 
         .Z(n11_adj_3724)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i2_2_lut_3_lut_adj_208.init = 16'h4040;
    LUT4 i2_2_lut_3_lut_adj_209 (.A(\operand_w[1] ), .B(size_w[0]), .C(data_w[29]), 
         .Z(n11_adj_3725)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i2_2_lut_3_lut_adj_209.init = 16'h4040;
    LUT4 i2_2_lut_3_lut_adj_210 (.A(\operand_w[1] ), .B(size_w[0]), .C(data_w[30]), 
         .Z(n11_adj_3726)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i2_2_lut_3_lut_adj_210.init = 16'h4040;
    LUT4 i1_2_lut_3_lut (.A(\operand_w[1] ), .B(size_w[0]), .C(data_w[31]), 
         .Z(n17)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_2_lut_3_lut.init = 16'h4040;
    FD1P3AX d_dat_o_i0_i28 (.D(store_data_m[28]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[28])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i28.GSR = "ENABLED";
    FD1P3AX d_dat_o_i0_i27 (.D(store_data_m[27]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[27])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i27.GSR = "ENABLED";
    FD1P3AX byte_enable_m_i0_i1 (.D(\byte_enable_x[1] ), .SP(w_clk_cpu_enable_972), 
            .CK(w_clk_cpu), .Q(byte_enable_m[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam byte_enable_m_i0_i1.GSR = "ENABLED";
    LUT4 i429_2_lut (.A(wb_load_complete_N_2129), .B(LM32D_CYC_O), .Z(w_clk_cpu_enable_438)) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(684[9] 733[12])
    defparam i429_2_lut.init = 16'h8888;
    LUT4 i56_3_lut (.A(n35), .B(data_w[16]), .C(size_w[1]), .Z(n32_adj_3727)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut (.A(sign_extend_w), .B(n41506), .C(size_w[1]), .Z(n27)) /* synthesis lut_function=(A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i56_3_lut_adj_211 (.A(n35), .B(data_w[17]), .C(size_w[1]), .Z(n32_adj_3728)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_211.init = 16'hcaca;
    FD1P3AX d_dat_o_i0_i26 (.D(store_data_m[26]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[26])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i26.GSR = "ENABLED";
    FD1P3AX d_dat_o_i0_i25 (.D(store_data_m[25]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[25])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i25.GSR = "ENABLED";
    FD1P3AX d_sel_o_i0_i3 (.D(byte_enable_m[3]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_SEL_O[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_sel_o_i0_i3.GSR = "ENABLED";
    LUT4 i56_3_lut_adj_212 (.A(n35), .B(data_w[18]), .C(size_w[1]), .Z(n32_adj_3729)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_212.init = 16'hcaca;
    LUT4 i56_3_lut_adj_213 (.A(n35), .B(data_w[19]), .C(size_w[1]), .Z(n32_adj_3730)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_213.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_3_lut (.A(size_w[0]), .B(data_w[14]), .C(\operand_w[1] ), 
         .Z(n36_adj_3731)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_2_lut_3_lut_3_lut.init = 16'hc4c4;
    FD1P3AX d_dat_o_i0_i24 (.D(store_data_m[24]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[24])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i24.GSR = "ENABLED";
    FD1P3AX d_dat_o_i0_i23 (.D(store_data_m[23]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[23])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i23.GSR = "ENABLED";
    FD1P3AX d_sel_o_i0_i2 (.D(byte_enable_m[2]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_SEL_O[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_sel_o_i0_i2.GSR = "ENABLED";
    LUT4 store_operand_x_5__bdd_4_lut (.A(store_operand_x[5]), .B(\size_x[1] ), 
         .C(store_operand_x[21]), .D(\condition_x[0] ), .Z(store_data_x[21])) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(((D)+!C)+!B)) */ ;
    defparam store_operand_x_5__bdd_4_lut.init = 16'h88e2;
    LUT4 i56_3_lut_adj_214 (.A(n35), .B(data_w[20]), .C(size_w[1]), .Z(n32_adj_3732)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_214.init = 16'hcaca;
    LUT4 i56_3_lut_adj_215 (.A(n35), .B(data_w[21]), .C(size_w[1]), .Z(n32_adj_3733)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_215.init = 16'hcaca;
    LUT4 i55_3_lut_adj_216 (.A(n32_adj_3733), .B(n27), .C(size_w[0]), 
         .Z(load_data_w[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_216.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut_adj_217 (.A(size_w[0]), .B(n31_adj_3734), .C(n25_adj_3711), 
         .D(size_w[1]), .Z(load_data_w[1])) /* synthesis lut_function=(A (C (D))+!A (B+(C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_217.init = 16'hf444;
    FD1P3AX d_dat_o_i0_i22 (.D(store_data_m[22]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[22])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i22.GSR = "ENABLED";
    FD1P3AX d_dat_o_i0_i21 (.D(store_data_m[21]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[21])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i21.GSR = "ENABLED";
    FD1P3AX d_sel_o_i0_i1 (.D(byte_enable_m[1]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_SEL_O[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_sel_o_i0_i1.GSR = "ENABLED";
    LUT4 i1_4_lut_4_lut_adj_218 (.A(size_w[0]), .B(n31_adj_3735), .C(n25_adj_3718), 
         .D(size_w[1]), .Z(load_data_w[3])) /* synthesis lut_function=(A (C (D))+!A (B+(C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_218.init = 16'hf444;
    LUT4 i1_4_lut_4_lut_adj_219 (.A(size_w[0]), .B(n31_adj_3736), .C(n25_adj_3715), 
         .D(size_w[1]), .Z(load_data_w[4])) /* synthesis lut_function=(A (C (D))+!A (B+(C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_219.init = 16'hf444;
    LUT4 i55_3_lut_adj_220 (.A(n32_adj_3732), .B(n27), .C(size_w[0]), 
         .Z(load_data_w[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_220.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_3_lut_adj_221 (.A(size_w[0]), .B(data_w[12]), .C(\operand_w[1] ), 
         .Z(n36_adj_3737)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_2_lut_3_lut_3_lut_adj_221.init = 16'hc4c4;
    LUT4 i1_2_lut_3_lut_3_lut_adj_222 (.A(size_w[0]), .B(data_w[8]), .C(\operand_w[1] ), 
         .Z(n36_adj_3738)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_2_lut_3_lut_3_lut_adj_222.init = 16'hc4c4;
    LUT4 i56_3_lut_adj_223 (.A(n35), .B(data_w[22]), .C(size_w[1]), .Z(n32_adj_3720)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_223.init = 16'hcaca;
    LUT4 i1_2_lut_3_lut_3_lut_adj_224 (.A(size_w[0]), .B(data_w[9]), .C(\operand_w[1] ), 
         .Z(n36_adj_3739)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_2_lut_3_lut_3_lut_adj_224.init = 16'hc4c4;
    LUT4 i56_3_lut_adj_225 (.A(n35), .B(data_w[23]), .C(size_w[1]), .Z(n32_adj_3719)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_225.init = 16'hcaca;
    LUT4 i56_3_lut_adj_226 (.A(n35), .B(data_w[24]), .C(size_w[1]), .Z(n32_adj_3709)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_226.init = 16'hcaca;
    FD1P3AX d_dat_o_i0_i20 (.D(store_data_m[20]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[20])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i20.GSR = "ENABLED";
    FD1P3AX d_dat_o_i0_i19 (.D(store_data_m[19]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[19])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i19.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_3_lut_adj_227 (.A(size_w[0]), .B(data_w[13]), .C(\operand_w[1] ), 
         .Z(n36_adj_3740)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_2_lut_3_lut_3_lut_adj_227.init = 16'hc4c4;
    LUT4 i1_2_lut_3_lut_3_lut_adj_228 (.A(size_w[0]), .B(data_w[11]), .C(\operand_w[1] ), 
         .Z(n36_adj_3741)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_2_lut_3_lut_3_lut_adj_228.init = 16'hc4c4;
    LUT4 i1_2_lut_2_lut (.A(size_w[0]), .B(n35), .Z(n33)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_2_lut_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_3_lut_3_lut_adj_229 (.A(size_w[0]), .B(data_w[10]), .C(\operand_w[1] ), 
         .Z(n36_adj_3742)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_2_lut_3_lut_3_lut_adj_229.init = 16'hc4c4;
    LUT4 i48_2_lut_3_lut_3_lut (.A(size_w[0]), .B(data_w[15]), .C(\operand_w[1] ), 
         .Z(n33_adj_3743)) /* synthesis lut_function=(A (B (C))+!A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i48_2_lut_3_lut_3_lut.init = 16'hc4c4;
    LUT4 i55_3_lut_adj_230 (.A(n32_adj_3730), .B(n27), .C(size_w[0]), 
         .Z(load_data_w[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_230.init = 16'hcaca;
    LUT4 i1_4_lut_4_lut_adj_231 (.A(size_w[0]), .B(n31_adj_3744), .C(n25_adj_3714), 
         .D(size_w[1]), .Z(load_data_w[5])) /* synthesis lut_function=(A (C (D))+!A (B+(C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_231.init = 16'hf444;
    FD1P3AX d_dat_o_i0_i18 (.D(store_data_m[18]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[18])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i18.GSR = "ENABLED";
    FD1P3AX d_dat_o_i0_i17 (.D(store_data_m[17]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[17])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i17.GSR = "ENABLED";
    LUT4 i1_4_lut_4_lut_adj_232 (.A(size_w[0]), .B(n31_adj_3707), .C(n25_adj_3713), 
         .D(size_w[1]), .Z(load_data_w[6])) /* synthesis lut_function=(A (C (D))+!A (B+(C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_232.init = 16'hf444;
    LUT4 i1_4_lut_4_lut_adj_233 (.A(size_w[0]), .B(n31), .C(n36), .D(size_w[1]), 
         .Z(load_data_w[7])) /* synthesis lut_function=(A (C (D))+!A (B+(C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_233.init = 16'hf444;
    LUT4 i1_4_lut_4_lut_adj_234 (.A(size_w[0]), .B(n31_adj_3745), .C(n25_adj_3716), 
         .D(size_w[1]), .Z(load_data_w[0])) /* synthesis lut_function=(A (C (D))+!A (B+(C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_234.init = 16'hf444;
    LUT4 i1_4_lut_4_lut_adj_235 (.A(size_w[0]), .B(n31_adj_3746), .C(n25), 
         .D(size_w[1]), .Z(load_data_w[2])) /* synthesis lut_function=(A (C (D))+!A (B+(C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_235.init = 16'hf444;
    FD1P3IX store_data_m_i0_i0 (.D(store_operand_x[0]), .SP(w_clk_cpu_enable_972), 
            .CD(n26122), .CK(w_clk_cpu), .Q(store_data_m[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i0.GSR = "ENABLED";
    LUT4 i55_3_lut_adj_236 (.A(n32_adj_3729), .B(n27), .C(size_w[0]), 
         .Z(load_data_w[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_236.init = 16'hcaca;
    FD1P3AX d_dat_o_i0_i16 (.D(store_data_m[16]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[16])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i16.GSR = "ENABLED";
    FD1P3AX d_dat_o_i0_i15 (.D(store_data_m[15]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[15])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i15.GSR = "ENABLED";
    FD1P3AX d_dat_o_i0_i14 (.D(store_data_m[14]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[14])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i14.GSR = "ENABLED";
    FD1P3AX d_dat_o_i0_i13 (.D(store_data_m[13]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[13])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i13.GSR = "ENABLED";
    LUT4 i55_3_lut_adj_237 (.A(n32_adj_3728), .B(n27), .C(size_w[0]), 
         .Z(load_data_w[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_237.init = 16'hcaca;
    FD1P3AX size_m_i0_i1 (.D(\size_x[1] ), .SP(w_clk_cpu_enable_711), .CK(w_clk_cpu), 
            .Q(size_m[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam size_m_i0_i1.GSR = "ENABLED";
    FD1P3AX d_dat_o_i0_i12 (.D(store_data_m[12]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[12])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i12.GSR = "ENABLED";
    FD1P3AX d_dat_o_i0_i11 (.D(store_data_m[11]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[11])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i11.GSR = "ENABLED";
    LUT4 i56_3_lut_adj_238 (.A(n35), .B(data_w[25]), .C(size_w[1]), .Z(n32_adj_3705)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_238.init = 16'hcaca;
    LUT4 store_operand_x_3__bdd_4_lut (.A(store_operand_x[3]), .B(\size_x[1] ), 
         .C(store_operand_x[19]), .D(\condition_x[0] ), .Z(store_data_x[19])) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(((D)+!C)+!B)) */ ;
    defparam store_operand_x_3__bdd_4_lut.init = 16'h88e2;
    LUT4 i56_3_lut_adj_239 (.A(n35), .B(data_w[26]), .C(size_w[1]), .Z(n32_adj_3704)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_239.init = 16'hcaca;
    FD1P3AX d_dat_o_i0_i10 (.D(store_data_m[10]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[10])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i10.GSR = "ENABLED";
    FD1P3AX d_dat_o_i0_i9 (.D(store_data_m[9]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[9])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i9.GSR = "ENABLED";
    LUT4 i56_3_lut_adj_240 (.A(n35), .B(data_w[27]), .C(size_w[1]), .Z(n32_adj_3703)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_240.init = 16'hcaca;
    LUT4 store_operand_x_2__bdd_4_lut (.A(store_operand_x[2]), .B(\size_x[1] ), 
         .C(store_operand_x[18]), .D(\condition_x[0] ), .Z(store_data_x[18])) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(((D)+!C)+!B)) */ ;
    defparam store_operand_x_2__bdd_4_lut.init = 16'h88e2;
    FD1P3AX d_dat_o_i0_i8 (.D(store_data_m[8]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[8])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i8.GSR = "ENABLED";
    FD1P3AX d_dat_o_i0_i7 (.D(store_data_m[7]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[7])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i7.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(stall_wb_load_N_2112), .B(n42746), .C(n46), .D(n4), 
         .Z(w_clk_cpu_enable_979)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;
    defparam i2_4_lut.init = 16'hefee;
    FD1P3AX d_dat_o_i0_i6 (.D(store_data_m[6]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[6])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i6.GSR = "ENABLED";
    FD1P3AX d_dat_o_i0_i5 (.D(store_data_m[5]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[5])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i5.GSR = "ENABLED";
    LUT4 i56_3_lut_adj_241 (.A(n35), .B(data_w[28]), .C(size_w[1]), .Z(n32_adj_3702)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_241.init = 16'hcaca;
    LUT4 i56_3_lut_adj_242 (.A(n35), .B(data_w[29]), .C(size_w[1]), .Z(n32)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_242.init = 16'hcaca;
    FD1P3AX d_dat_o_i0_i4 (.D(store_data_m[4]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i4.GSR = "ENABLED";
    FD1P3AX d_dat_o_i0_i3 (.D(store_data_m[3]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i3.GSR = "ENABLED";
    LUT4 i56_3_lut_adj_243 (.A(n35), .B(data_w[30]), .C(size_w[1]), .Z(n32_adj_3747)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_243.init = 16'hcaca;
    LUT4 store_operand_x_4__bdd_4_lut (.A(store_operand_x[4]), .B(\size_x[1] ), 
         .C(store_operand_x[20]), .D(\condition_x[0] ), .Z(store_data_x[20])) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(((D)+!C)+!B)) */ ;
    defparam store_operand_x_4__bdd_4_lut.init = 16'h88e2;
    FD1P3AX d_dat_o_i0_i2 (.D(store_data_m[2]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i2.GSR = "ENABLED";
    FD1P3AX d_dat_o_i0_i1 (.D(store_data_m[1]), .SP(w_clk_cpu_enable_623), 
            .CK(w_clk_cpu), .Q(LM32D_DAT_O[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_dat_o_i0_i1.GSR = "ENABLED";
    FD1S3AX data_w_i31 (.D(data_m[31]), .CK(w_clk_cpu), .Q(data_w[31])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i31.GSR = "ENABLED";
    FD1S3AX data_w_i30 (.D(data_m[30]), .CK(w_clk_cpu), .Q(data_w[30])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i30.GSR = "ENABLED";
    FD1S3AX data_w_i29 (.D(data_m[29]), .CK(w_clk_cpu), .Q(data_w[29])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i29.GSR = "ENABLED";
    FD1S3AX data_w_i28 (.D(data_m[28]), .CK(w_clk_cpu), .Q(data_w[28])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i28.GSR = "ENABLED";
    FD1S3AX data_w_i27 (.D(data_m[27]), .CK(w_clk_cpu), .Q(data_w[27])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i27.GSR = "ENABLED";
    LUT4 i56_3_lut_adj_244 (.A(n35), .B(data_w[31]), .C(size_w[1]), .Z(n32_adj_3748)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i56_3_lut_adj_244.init = 16'hcaca;
    PFUMX i52_adj_245 (.BLUT(n23_adj_3749), .ALUT(n28_adj_3750), .C0(\operand_w[1] ), 
          .Z(n31_adj_3745));
    FD1S3AX data_w_i26 (.D(data_m[26]), .CK(w_clk_cpu), .Q(data_w[26])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i26.GSR = "ENABLED";
    FD1S3AX data_w_i25 (.D(data_m[25]), .CK(w_clk_cpu), .Q(data_w[25])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i25.GSR = "ENABLED";
    FD1S3AX data_w_i24 (.D(data_m[24]), .CK(w_clk_cpu), .Q(data_w[24])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i24.GSR = "ENABLED";
    FD1S3AX data_w_i23 (.D(data_m[23]), .CK(w_clk_cpu), .Q(data_w[23])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i23.GSR = "ENABLED";
    PFUMX i52_adj_246 (.BLUT(n23_adj_3751), .ALUT(n28_adj_3752), .C0(\operand_w[1] ), 
          .Z(n31_adj_3735));
    PFUMX i52_adj_247 (.BLUT(n23_adj_3753), .ALUT(n28_adj_3754), .C0(\operand_w[1] ), 
          .Z(n31_adj_3734));
    LUT4 i33847_3_lut_rep_418 (.A(data_w[23]), .B(data_w[7]), .C(\operand_w[1] ), 
         .Z(n41505)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(527[22:31])
    defparam i33847_3_lut_rep_418.init = 16'hcaca;
    LUT4 i31_4_lut_4_lut_4_lut (.A(data_w[23]), .B(data_w[7]), .C(\operand_w[1] ), 
         .D(size_w[1]), .Z(n28)) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(527[22:31])
    defparam i31_4_lut_4_lut_4_lut.init = 16'hc0ca;
    FD1S3AX data_w_i22 (.D(data_m[22]), .CK(w_clk_cpu), .Q(data_w[22])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i22.GSR = "ENABLED";
    FD1S3AX data_w_i21 (.D(data_m[21]), .CK(w_clk_cpu), .Q(data_w[21])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i21.GSR = "ENABLED";
    LUT4 i33842_3_lut_rep_419 (.A(data_w[31]), .B(data_w[15]), .C(\operand_w[1] ), 
         .Z(n41506)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(527[22:31])
    defparam i33842_3_lut_rep_419.init = 16'hcaca;
    LUT4 i1_2_lut_2_lut_4_lut (.A(data_w[31]), .B(data_w[15]), .C(\operand_w[1] ), 
         .D(size_w[1]), .Z(n30)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(527[22:31])
    defparam i1_2_lut_2_lut_4_lut.init = 16'h00ca;
    FD1S3AX data_w_i20 (.D(data_m[20]), .CK(w_clk_cpu), .Q(data_w[20])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i20.GSR = "ENABLED";
    FD1S3AX data_w_i19 (.D(data_m[19]), .CK(w_clk_cpu), .Q(data_w[19])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i19.GSR = "ENABLED";
    PFUMX i52_adj_248 (.BLUT(n23_adj_3755), .ALUT(n28_adj_3756), .C0(\operand_w[1] ), 
          .Z(n31_adj_3736));
    LUT4 size_x_1__I_0_153_Mux_8_i3_3_lut_4_lut (.A(store_operand_x[0]), .B(\condition_x[0] ), 
         .C(\size_x[1] ), .D(store_operand_x[8]), .Z(store_data_x[8])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_153_Mux_8_i3_3_lut_4_lut.init = 16'hf202;
    LUT4 size_x_1__I_0_153_Mux_24_i3_3_lut_4_lut (.A(store_operand_x[0]), 
         .B(\condition_x[0] ), .C(\size_x[1] ), .D(n2_adj_3717), .Z(store_data_x[24])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_153_Mux_24_i3_3_lut_4_lut.init = 16'hf202;
    FD1S3AX data_w_i18 (.D(data_m[18]), .CK(w_clk_cpu), .Q(data_w[18])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i18.GSR = "ENABLED";
    FD1S3AX data_w_i17 (.D(data_m[17]), .CK(w_clk_cpu), .Q(data_w[17])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i17.GSR = "ENABLED";
    LUT4 i21704_3_lut (.A(wb_load_complete_N_2129), .B(n41428), .C(LM32D_CYC_O), 
         .Z(w_clk_cpu_enable_27)) /* synthesis lut_function=(A ((C)+!B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam i21704_3_lut.init = 16'ha2a2;
    FD1S3AX data_w_i16 (.D(data_m[16]), .CK(w_clk_cpu), .Q(data_w[16])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i16.GSR = "ENABLED";
    FD1S3AX data_w_i15 (.D(data_m[15]), .CK(w_clk_cpu), .Q(data_w[15])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i15.GSR = "ENABLED";
    LUT4 d_we_o_I_0_1_lut (.A(LM32D_WE_O), .Z(d_we_o_N_2124)) /* synthesis lut_function=(!(A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(676[40:47])
    defparam d_we_o_I_0_1_lut.init = 16'h5555;
    PFUMX i52_adj_249 (.BLUT(n23_adj_3757), .ALUT(n28_adj_3758), .C0(\operand_w[1] ), 
          .Z(n31_adj_3746));
    LUT4 store_operand_x_7__bdd_4_lut (.A(store_operand_x[7]), .B(\size_x[1] ), 
         .C(store_operand_x[23]), .D(\condition_x[0] ), .Z(store_data_x[23])) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(((D)+!C)+!B)) */ ;
    defparam store_operand_x_7__bdd_4_lut.init = 16'h88e2;
    LUT4 size_x_1__I_0_153_Mux_9_i3_3_lut_4_lut (.A(store_operand_x[1]), .B(\condition_x[0] ), 
         .C(\size_x[1] ), .D(store_operand_x[9]), .Z(store_data_x[9])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_153_Mux_9_i3_3_lut_4_lut.init = 16'hf202;
    FD1S3AX data_w_i14 (.D(data_m[14]), .CK(w_clk_cpu), .Q(data_w[14])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i14.GSR = "ENABLED";
    LUT4 size_x_1__I_0_153_Mux_25_i3_3_lut_4_lut (.A(store_operand_x[1]), 
         .B(\condition_x[0] ), .C(\size_x[1] ), .D(n2_adj_3712), .Z(store_data_x[25])) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(449[5] 454[12])
    defparam size_x_1__I_0_153_Mux_25_i3_3_lut_4_lut.init = 16'hf202;
    PFUMX i52_adj_250 (.BLUT(n23_adj_3759), .ALUT(n28_adj_3760), .C0(\operand_w[1] ), 
          .Z(n31_adj_3744));
    FD1P3IX store_data_m_i0_i2 (.D(store_operand_x[2]), .SP(w_clk_cpu_enable_972), 
            .CD(n26122), .CK(w_clk_cpu), .Q(store_data_m[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i2.GSR = "ENABLED";
    FD1S3AX data_w_i13 (.D(data_m[13]), .CK(w_clk_cpu), .Q(data_w[13])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i13.GSR = "ENABLED";
    FD1S3AX data_w_i12 (.D(data_m[12]), .CK(w_clk_cpu), .Q(data_w[12])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i12.GSR = "ENABLED";
    FD1S3AX data_w_i11 (.D(data_m[11]), .CK(w_clk_cpu), .Q(data_w[11])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i11.GSR = "ENABLED";
    FD1S3AX data_w_i10 (.D(data_m[10]), .CK(w_clk_cpu), .Q(data_w[10])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i10.GSR = "ENABLED";
    LUT4 i38022_3_lut_4_lut (.A(n41491), .B(\adder_result_x[1] ), .C(n32389), 
         .D(\adder_result_x[0] ), .Z(byte_enable_x_c[3])) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C (D))))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(464[5:29])
    defparam i38022_3_lut_4_lut.init = 16'h0f1f;
    LUT4 i1_3_lut_4_lut (.A(n41491), .B(\adder_result_x[1] ), .C(n32389), 
         .D(\adder_result_x[0] ), .Z(byte_enable_x_c[2])) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !((D)+!C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(464[5:29])
    defparam i1_3_lut_4_lut.init = 16'h1f0f;
    FD1S3AX data_w_i9 (.D(data_m[9]), .CK(w_clk_cpu), .Q(data_w[9])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i9.GSR = "ENABLED";
    FD1S3AX data_w_i8 (.D(data_m[8]), .CK(w_clk_cpu), .Q(data_w[8])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i8.GSR = "ENABLED";
    LUT4 i55_3_lut_adj_251 (.A(n32_adj_3748), .B(n27), .C(size_w[0]), 
         .Z(load_data_w[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_251.init = 16'hcaca;
    LUT4 i55_3_lut_adj_252 (.A(n32_adj_3747), .B(n27), .C(size_w[0]), 
         .Z(load_data_w[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_252.init = 16'hcaca;
    LUT4 i55_3_lut_adj_253 (.A(n32_adj_3727), .B(n27), .C(size_w[0]), 
         .Z(load_data_w[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i55_3_lut_adj_253.init = 16'hcaca;
    FD1P3AX d_adr_o_i0_i31 (.D(operand_m[31]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[31])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i31.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i30 (.D(operand_m[30]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[30])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i30.GSR = "ENABLED";
    FD1S3AX data_w_i7 (.D(data_m[7]), .CK(w_clk_cpu), .Q(data_w[7])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i7.GSR = "ENABLED";
    LUT4 i33861_4_lut (.A(n33), .B(n33_adj_3743), .C(size_w[1]), .D(n17), 
         .Z(load_data_w[15])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(240[22:28])
    defparam i33861_4_lut.init = 16'hfaca;
    LUT4 store_operand_x_6__bdd_4_lut (.A(store_operand_x[6]), .B(\size_x[1] ), 
         .C(store_operand_x[22]), .D(\condition_x[0] ), .Z(store_data_x[22])) /* synthesis lut_function=(A (B (C+(D))+!B !(D))+!A !(((D)+!C)+!B)) */ ;
    defparam store_operand_x_6__bdd_4_lut.init = 16'h88e2;
    FD1P3AX d_adr_o_i0_i29 (.D(operand_m[29]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[29])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i29.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i28 (.D(operand_m[28]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[28])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i28.GSR = "ENABLED";
    FD1S3AX data_w_i6 (.D(data_m[6]), .CK(w_clk_cpu), .Q(data_w[6])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i6.GSR = "ENABLED";
    FD1P3IX store_data_m_i0_i3 (.D(store_operand_x[3]), .SP(w_clk_cpu_enable_972), 
            .CD(n26122), .CK(w_clk_cpu), .Q(store_data_m[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i3.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i27 (.D(operand_m[27]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[27])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i27.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i26 (.D(operand_m[26]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[26])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i26.GSR = "ENABLED";
    FD1S3AX data_w_i5 (.D(data_m[5]), .CK(w_clk_cpu), .Q(data_w[5])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i5.GSR = "ENABLED";
    LUT4 i53_4_lut (.A(n33), .B(n11_adj_3726), .C(size_w[1]), .D(n36_adj_3731), 
         .Z(load_data_w[14])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut.init = 16'hfaca;
    FD1P3AX d_adr_o_i0_i25 (.D(operand_m[25]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[25])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i25.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i24 (.D(operand_m[24]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[24])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i24.GSR = "ENABLED";
    FD1S3AX data_w_i4 (.D(data_m[4]), .CK(w_clk_cpu), .Q(data_w[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i4.GSR = "ENABLED";
    LUT4 i53_4_lut_adj_254 (.A(n33), .B(n11_adj_3725), .C(size_w[1]), 
         .D(n36_adj_3740), .Z(load_data_w[13])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut_adj_254.init = 16'hfaca;
    FD1P3IX store_data_m_i0_i4 (.D(store_operand_x[4]), .SP(w_clk_cpu_enable_972), 
            .CD(n26122), .CK(w_clk_cpu), .Q(store_data_m[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i4.GSR = "ENABLED";
    LUT4 i53_4_lut_adj_255 (.A(n33), .B(n11_adj_3724), .C(size_w[1]), 
         .D(n36_adj_3737), .Z(load_data_w[12])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut_adj_255.init = 16'hfaca;
    FD1P3AX d_adr_o_i0_i23 (.D(operand_m[23]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[23])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i23.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i22 (.D(operand_m[22]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[22])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i22.GSR = "ENABLED";
    FD1S3AX data_w_i3 (.D(data_m[3]), .CK(w_clk_cpu), .Q(data_w[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i3.GSR = "ENABLED";
    LUT4 i53_4_lut_adj_256 (.A(n33), .B(n11_adj_3722), .C(size_w[1]), 
         .D(n36_adj_3741), .Z(load_data_w[11])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut_adj_256.init = 16'hfaca;
    FD1P3AX d_adr_o_i0_i21 (.D(operand_m[21]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[21])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i21.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i20 (.D(operand_m[20]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[20])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i20.GSR = "ENABLED";
    FD1S3AX data_w_i2 (.D(data_m[2]), .CK(w_clk_cpu), .Q(data_w[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i2.GSR = "ENABLED";
    FD1P3AX wb_select_m_141 (.D(n42726), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(wb_select_m));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam wb_select_m_141.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i19 (.D(operand_m[19]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[19])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i19.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i18 (.D(operand_m[18]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[18])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i18.GSR = "ENABLED";
    FD1S3AX data_w_i1 (.D(data_m[1]), .CK(w_clk_cpu), .Q(data_w[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam data_w_i1.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i17 (.D(operand_m[17]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[17])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i17.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i16 (.D(operand_m[16]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[16])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i16.GSR = "ENABLED";
    FD1S3AX size_w_i1 (.D(size_m[1]), .CK(w_clk_cpu), .Q(size_w[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(800[5] 804[8])
    defparam size_w_i1.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i15 (.D(operand_m[15]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[15])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i15.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i14 (.D(operand_m[14]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[14])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i14.GSR = "ENABLED";
    FD1P3AX store_data_m_i0_i31 (.D(\store_data_x[31] ), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(store_data_m[31])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i31.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i13 (.D(operand_m[13]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[13])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i13.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i12 (.D(operand_m[12]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[12])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i12.GSR = "ENABLED";
    FD1P3AX store_data_m_i0_i30 (.D(\store_data_x[30] ), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(store_data_m[30])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i30.GSR = "ENABLED";
    FD1P3AX sign_extend_m_137 (.D(sign_extend_x), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(sign_extend_m));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam sign_extend_m_137.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i11 (.D(operand_m[11]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[11])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i11.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i10 (.D(operand_m[10]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[10])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i10.GSR = "ENABLED";
    FD1P3AX store_data_m_i0_i29 (.D(store_data_x[29]), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(store_data_m[29])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i29.GSR = "ENABLED";
    LUT4 i53_4_lut_adj_257 (.A(n33), .B(n11_adj_3723), .C(size_w[1]), 
         .D(n36_adj_3742), .Z(load_data_w[10])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut_adj_257.init = 16'hfaca;
    FD1P3AX d_adr_o_i0_i9 (.D(operand_m[9]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[9])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i9.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i8 (.D(operand_m[8]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[8])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i8.GSR = "ENABLED";
    FD1P3AX store_data_m_i0_i28 (.D(store_data_x[28]), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(store_data_m[28])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i28.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i7 (.D(operand_m[7]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[7])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i7.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i6 (.D(operand_m[6]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[6])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i6.GSR = "ENABLED";
    FD1P3AX store_data_m_i0_i27 (.D(store_data_x[27]), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(store_data_m[27])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i27.GSR = "ENABLED";
    LUT4 i53_4_lut_adj_258 (.A(n33), .B(n11_adj_3721), .C(size_w[1]), 
         .D(n36_adj_3739), .Z(load_data_w[9])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut_adj_258.init = 16'hfaca;
    FD1P3AX d_adr_o_i0_i5 (.D(operand_m[5]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[5])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i5.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i4 (.D(operand_m[4]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i4.GSR = "ENABLED";
    FD1P3AX store_data_m_i0_i26 (.D(store_data_x[26]), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(store_data_m[26])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i26.GSR = "ENABLED";
    FD1P3IX store_data_m_i0_i5 (.D(store_operand_x[5]), .SP(w_clk_cpu_enable_972), 
            .CD(n26122), .CK(w_clk_cpu), .Q(store_data_m[5])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i5.GSR = "ENABLED";
    LUT4 i1_3_lut (.A(\condition_x[0] ), .B(\size_x[1] ), .C(\adder_result_x[1] ), 
         .Z(n32389)) /* synthesis lut_function=(A ((C)+!B)+!A !(B)) */ ;
    defparam i1_3_lut.init = 16'hb3b3;
    FD1P3AX d_adr_o_i0_i3 (.D(operand_m[3]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i3.GSR = "ENABLED";
    FD1P3AX d_adr_o_i0_i2 (.D(operand_m[2]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i2.GSR = "ENABLED";
    FD1P3AX store_data_m_i0_i25 (.D(store_data_x[25]), .SP(w_clk_cpu_enable_878), 
            .CK(w_clk_cpu), .Q(store_data_m[25])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i25.GSR = "ENABLED";
    LUT4 i53_4_lut_adj_259 (.A(n33), .B(n11), .C(size_w[1]), .D(n36_adj_3738), 
         .Z(load_data_w[8])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut_adj_259.init = 16'hfaca;
    FD1P3AX d_adr_o_i0_i1 (.D(operand_m[1]), .SP(w_clk_cpu_enable_886), 
            .CK(w_clk_cpu), .Q(LM32D_ADR_O[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam d_adr_o_i0_i1.GSR = "ENABLED";
    FD1P3AX store_data_m_i0_i24 (.D(store_data_x[24]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(store_data_m[24])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i24.GSR = "ENABLED";
    FD1P3AX store_data_m_i0_i23 (.D(store_data_x[23]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(store_data_m[23])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i23.GSR = "ENABLED";
    LUT4 i1_4_lut_4_lut_adj_260 (.A(size_w[1]), .B(\operand_w[0] ), .C(data_w[18]), 
         .D(data_w[26]), .Z(n23_adj_3757)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_260.init = 16'h5140;
    FD1P3AX store_data_m_i0_i22 (.D(store_data_x[22]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(store_data_m[22])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i22.GSR = "ENABLED";
    LUT4 i53_4_lut_4_lut (.A(size_w[1]), .B(data_w[14]), .C(\operand_w[0] ), 
         .D(data_w[6]), .Z(n28_adj_3706)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut_4_lut.init = 16'hf404;
    LUT4 i1_4_lut_4_lut_adj_261 (.A(size_w[1]), .B(\operand_w[0] ), .C(data_w[17]), 
         .D(data_w[25]), .Z(n23_adj_3753)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_261.init = 16'h5140;
    LUT4 i1_4_lut_4_lut_adj_262 (.A(size_w[1]), .B(\operand_w[0] ), .C(data_w[20]), 
         .D(data_w[28]), .Z(n23_adj_3755)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_262.init = 16'h5140;
    LUT4 i1_4_lut_4_lut_adj_263 (.A(size_w[1]), .B(\operand_w[0] ), .C(data_w[21]), 
         .D(data_w[29]), .Z(n23_adj_3759)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_263.init = 16'h5140;
    LUT4 i53_4_lut_4_lut_adj_264 (.A(size_w[1]), .B(data_w[8]), .C(\operand_w[0] ), 
         .D(data_w[0]), .Z(n28_adj_3750)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut_4_lut_adj_264.init = 16'hf404;
    LUT4 i53_4_lut_4_lut_adj_265 (.A(size_w[1]), .B(data_w[10]), .C(\operand_w[0] ), 
         .D(data_w[2]), .Z(n28_adj_3758)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut_4_lut_adj_265.init = 16'hf404;
    LUT4 i1_4_lut_4_lut_adj_266 (.A(size_w[1]), .B(\operand_w[0] ), .C(data_w[16]), 
         .D(data_w[24]), .Z(n23_adj_3749)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_266.init = 16'h5140;
    LUT4 i53_4_lut_4_lut_adj_267 (.A(size_w[1]), .B(data_w[12]), .C(\operand_w[0] ), 
         .D(data_w[4]), .Z(n28_adj_3756)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut_4_lut_adj_267.init = 16'hf404;
    FD1P3AX store_data_m_i0_i21 (.D(store_data_x[21]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(store_data_m[21])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i21.GSR = "ENABLED";
    LUT4 i53_4_lut_4_lut_adj_268 (.A(size_w[1]), .B(data_w[9]), .C(\operand_w[0] ), 
         .D(data_w[1]), .Z(n28_adj_3754)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut_4_lut_adj_268.init = 16'hf404;
    LUT4 i53_4_lut_4_lut_adj_269 (.A(size_w[1]), .B(data_w[13]), .C(\operand_w[0] ), 
         .D(data_w[5]), .Z(n28_adj_3760)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut_4_lut_adj_269.init = 16'hf404;
    LUT4 i1_4_lut_4_lut_adj_270 (.A(size_w[1]), .B(\operand_w[0] ), .C(data_w[19]), 
         .D(data_w[27]), .Z(n23_adj_3751)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_270.init = 16'h5140;
    LUT4 i53_4_lut_4_lut_adj_271 (.A(size_w[1]), .B(data_w[11]), .C(\operand_w[0] ), 
         .D(data_w[3]), .Z(n28_adj_3752)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i53_4_lut_4_lut_adj_271.init = 16'hf404;
    LUT4 i1_4_lut_4_lut_adj_272 (.A(size_w[1]), .B(\operand_w[0] ), .C(data_w[22]), 
         .D(data_w[30]), .Z(n23)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(574[5] 583[12])
    defparam i1_4_lut_4_lut_adj_272.init = 16'h5140;
    FD1P3AX store_data_m_i0_i20 (.D(store_data_x[20]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(store_data_m[20])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i20.GSR = "ENABLED";
    FD1P3AX store_data_m_i0_i19 (.D(store_data_x[19]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(store_data_m[19])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i19.GSR = "ENABLED";
    FD1P3AX store_data_m_i0_i18 (.D(store_data_x[18]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(store_data_m[18])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i18.GSR = "ENABLED";
    FD1P3AX store_data_m_i0_i17 (.D(store_data_x[17]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(store_data_m[17])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i17.GSR = "ENABLED";
    FD1P3AX store_data_m_i0_i16 (.D(store_data_x[16]), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(store_data_m[16])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i16.GSR = "ENABLED";
    FD1P3IX store_data_m_i0_i6 (.D(store_operand_x[6]), .SP(w_clk_cpu_enable_972), 
            .CD(n26122), .CK(w_clk_cpu), .Q(store_data_m[6])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i6.GSR = "ENABLED";
    FD1P3IX store_data_m_i0_i7 (.D(store_operand_x[7]), .SP(w_clk_cpu_enable_972), 
            .CD(n26122), .CK(w_clk_cpu), .Q(store_data_m[7])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i7.GSR = "ENABLED";
    FD1P3AX store_data_m_i0_i15 (.D(\store_data_x[15] ), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(store_data_m[15])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i15.GSR = "ENABLED";
    FD1P3IX stall_wb_load_136 (.D(stall_wb_load_N_2112), .SP(w_clk_cpu_enable_979), 
            .CD(exception_m), .CK(w_clk_cpu), .Q(stall_wb_load));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(643[5] 743[8])
    defparam stall_wb_load_136.GSR = "ENABLED";
    FD1P3AX store_data_m_i0_i14 (.D(\store_data_x[14] ), .SP(w_clk_cpu_enable_985), 
            .CK(w_clk_cpu), .Q(store_data_m[14])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=984, LSE_RLINE=1043 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_load_store_unit.v(769[5] 787[8])
    defparam store_data_m_i0_i14.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module lm32_jtag
//

module lm32_jtag (jtag_reg_d, w_clk_cpu, GND_net, n41428, n39970, 
            branch_flushX_m_N_1116, cycles_5__N_2495, n42740, w_clk_cpu_enable_914, 
            n41391, load_x, n41395, stall_wb_load_N_2112, w_clk_cpu_enable_697, 
            n26126, csr_write_enable_x, n41357, LM32I_CYC_O, w_clk_cpu_enable_763, 
            branch_taken_m, w_clk_cpu_enable_638, w_clk_cpu_enable_984, 
            n41365, \csr_x[0] , n41444, n41457, eba_31__N_1101, \operand_1_x[0] , 
            n31712, deba_31__N_1120, jtag_break, reset_exception, \jrx_csr_read_data[0] , 
            jtag_reg_q, jtag_update_N_2932, \jtag_reg_addr_d[1] , \jtag_reg_addr_d[0] , 
            w_clk_cpu_enable_330, n42726, \jrx_csr_read_data[7] , \jrx_csr_read_data[6] , 
            \jrx_csr_read_data[5] , \jrx_csr_read_data[4] , \jrx_csr_read_data[3] , 
            \jrx_csr_read_data[2] , \jrx_csr_read_data[1] , w_clk_cpu_enable_865, 
            w_clk_cpu_enable_958, x_result_sel_csr_d, n22501, n41417, 
            n26142, w_clk_cpu_enable_983, jtag_reg_addr_q, n38725, jtag_reg_d_7__N_505, 
            \operand_1_x[7] , \operand_1_x[6] , \operand_1_x[5] , \operand_1_x[4] , 
            \operand_1_x[3] , \operand_1_x[2] , \operand_1_x[1] ) /* synthesis syn_module_defined=1 */ ;
    output [7:0]jtag_reg_d;
    input w_clk_cpu;
    input GND_net;
    input n41428;
    input n39970;
    input branch_flushX_m_N_1116;
    input cycles_5__N_2495;
    output n42740;
    output w_clk_cpu_enable_914;
    input n41391;
    input load_x;
    input n41395;
    output stall_wb_load_N_2112;
    input w_clk_cpu_enable_697;
    output n26126;
    input csr_write_enable_x;
    output n41357;
    input LM32I_CYC_O;
    output w_clk_cpu_enable_763;
    input branch_taken_m;
    output w_clk_cpu_enable_638;
    output w_clk_cpu_enable_984;
    input n41365;
    input \csr_x[0] ;
    input n41444;
    input n41457;
    output eba_31__N_1101;
    input \operand_1_x[0] ;
    input n31712;
    output deba_31__N_1120;
    output jtag_break;
    output reset_exception;
    output \jrx_csr_read_data[0] ;
    input [7:0]jtag_reg_q;
    input jtag_update_N_2932;
    output \jtag_reg_addr_d[1] ;
    output \jtag_reg_addr_d[0] ;
    input w_clk_cpu_enable_330;
    input n42726;
    output \jrx_csr_read_data[7] ;
    output \jrx_csr_read_data[6] ;
    output \jrx_csr_read_data[5] ;
    output \jrx_csr_read_data[4] ;
    output \jrx_csr_read_data[3] ;
    output \jrx_csr_read_data[2] ;
    output \jrx_csr_read_data[1] ;
    output w_clk_cpu_enable_865;
    output w_clk_cpu_enable_958;
    input x_result_sel_csr_d;
    output n22501;
    input n41417;
    output n26142;
    output w_clk_cpu_enable_983;
    input [2:0]jtag_reg_addr_q;
    input n38725;
    input jtag_reg_d_7__N_505;
    input \operand_1_x[7] ;
    input \operand_1_x[6] ;
    input \operand_1_x[5] ;
    input \operand_1_x[4] ;
    input \operand_1_x[3] ;
    input \operand_1_x[2] ;
    input \operand_1_x[1] ;
    
    wire w_clk_cpu /* synthesis SET_AS_NETWORK=w_clk_cpu, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(22[6:15])
    wire jtag_update_N_2932 /* synthesis is_inv_clock=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(203[14:23])
    
    wire w_clk_cpu_enable_872;
    wire [7:0]uart_tx_byte;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(212[28:40])
    
    wire w_clk_cpu_enable_769, rx_toggle_r, rx_toggle, rx_toggle_r_r, 
        rx_toggle_r_r_r, w_clk_cpu_enable_270, n41400, w_clk_cpu_enable_271, 
        n41399, jrx_csr_read_data_8__N_2865, rx_toggle_N_2930, w_clk_cpu_enable_275, 
        n24867, n41443, n40543, n41484, n41483, n25688, n38722, 
        n39169, n4, n10;
    
    FD1P3IX jtag_reg_d_i1 (.D(uart_tx_byte[1]), .SP(w_clk_cpu_enable_872), 
            .CD(GND_net), .CK(w_clk_cpu), .Q(jtag_reg_d[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam jtag_reg_d_i1.GSR = "ENABLED";
    FD1P3IX jtag_reg_d_i2 (.D(uart_tx_byte[2]), .SP(w_clk_cpu_enable_872), 
            .CD(GND_net), .CK(w_clk_cpu), .Q(jtag_reg_d[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam jtag_reg_d_i2.GSR = "ENABLED";
    FD1P3IX jtag_reg_d_i6 (.D(uart_tx_byte[6]), .SP(w_clk_cpu_enable_872), 
            .CD(GND_net), .CK(w_clk_cpu), .Q(jtag_reg_d[6])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam jtag_reg_d_i6.GSR = "ENABLED";
    LUT4 i37889_2_lut_rep_459 (.A(n41428), .B(n39970), .C(branch_flushX_m_N_1116), 
         .D(cycles_5__N_2495), .Z(n42740)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2421[13:30])
    defparam i37889_2_lut_rep_459.init = 16'h4440;
    LUT4 i37889_2_lut_rep_460 (.A(n41428), .B(n39970), .C(branch_flushX_m_N_1116), 
         .D(cycles_5__N_2495), .Z(w_clk_cpu_enable_914)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2421[13:30])
    defparam i37889_2_lut_rep_460.init = 16'h4440;
    LUT4 i1_3_lut_4_lut_4_lut (.A(n41428), .B(n41391), .C(load_x), .D(n41395), 
         .Z(stall_wb_load_N_2112)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2421[13:30])
    defparam i1_3_lut_4_lut_4_lut.init = 16'h4000;
    LUT4 i23485_2_lut_2_lut_3_lut_4_lut_4_lut (.A(n41428), .B(n39970), .C(w_clk_cpu_enable_697), 
         .D(n41395), .Z(n26126)) /* synthesis lut_function=(A (C)+!A !(B ((D)+!C)+!B !(C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2421[13:30])
    defparam i23485_2_lut_2_lut_3_lut_4_lut_4_lut.init = 16'hb0f0;
    LUT4 i1_2_lut_rep_270_3_lut_4_lut_4_lut (.A(n41428), .B(csr_write_enable_x), 
         .C(n41391), .D(n41395), .Z(n41357)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2421[13:30])
    defparam i1_2_lut_rep_270_3_lut_4_lut_4_lut.init = 16'h4000;
    LUT4 i37837_2_lut_3_lut_4_lut_4_lut (.A(n41428), .B(n39970), .C(LM32I_CYC_O), 
         .D(n41395), .Z(w_clk_cpu_enable_763)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2421[13:30])
    defparam i37837_2_lut_3_lut_4_lut_4_lut.init = 16'h0400;
    FD1P3IX jtag_reg_d_i7 (.D(uart_tx_byte[7]), .SP(w_clk_cpu_enable_872), 
            .CD(GND_net), .CK(w_clk_cpu), .Q(jtag_reg_d[7])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam jtag_reg_d_i7.GSR = "ENABLED";
    LUT4 i19862_2_lut_3_lut_4_lut_4_lut (.A(n41428), .B(n39970), .C(branch_taken_m), 
         .D(n41395), .Z(w_clk_cpu_enable_638)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2421[13:30])
    defparam i19862_2_lut_3_lut_4_lut_4_lut.init = 16'hf4f0;
    LUT4 i37893_2_lut_rep_290_3_lut_4_lut_3_lut (.A(n41428), .B(cycles_5__N_2495), 
         .C(branch_flushX_m_N_1116), .Z(w_clk_cpu_enable_984)) /* synthesis lut_function=(!(A+!(B+(C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2421[13:30])
    defparam i37893_2_lut_rep_290_3_lut_4_lut_3_lut.init = 16'h5454;
    LUT4 i2_3_lut_4_lut (.A(n41365), .B(w_clk_cpu_enable_984), .C(\csr_x[0] ), 
         .D(n41444), .Z(w_clk_cpu_enable_769)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(341[18:68])
    defparam i2_3_lut_4_lut.init = 16'h0800;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n41365), .B(w_clk_cpu_enable_984), .C(n41457), 
         .D(\csr_x[0] ), .Z(eba_31__N_1101)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(341[18:68])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h8000;
    FD1P3AX uart_tx_byte_i0_i0 (.D(\operand_1_x[0] ), .SP(w_clk_cpu_enable_769), 
            .CK(w_clk_cpu), .Q(uart_tx_byte[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_tx_byte_i0_i0.GSR = "ENABLED";
    FD1S3AX rx_toggle_r_82 (.D(rx_toggle), .CK(w_clk_cpu), .Q(rx_toggle_r)) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(301[4] 305[7])
    defparam rx_toggle_r_82.GSR = "ENABLED";
    FD1S3AX rx_toggle_r_r_83 (.D(rx_toggle_r), .CK(w_clk_cpu), .Q(rx_toggle_r_r)) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(301[4] 305[7])
    defparam rx_toggle_r_r_83.GSR = "ENABLED";
    FD1S3AX rx_toggle_r_r_r_84 (.D(rx_toggle_r_r), .CK(w_clk_cpu), .Q(rx_toggle_r_r_r)) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(301[4] 305[7])
    defparam rx_toggle_r_r_r_84.GSR = "ENABLED";
    FD1P3IX jtag_reg_d_i3 (.D(uart_tx_byte[3]), .SP(w_clk_cpu_enable_872), 
            .CD(GND_net), .CK(w_clk_cpu), .Q(jtag_reg_d[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam jtag_reg_d_i3.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut_adj_188 (.A(n41365), .B(w_clk_cpu_enable_984), 
         .C(n31712), .D(\csr_x[0] ), .Z(deba_31__N_1120)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(341[18:68])
    defparam i1_2_lut_3_lut_4_lut_adj_188.init = 16'h0800;
    FD1P3AX jtag_break_88 (.D(n41400), .SP(w_clk_cpu_enable_270), .CK(w_clk_cpu), 
            .Q(jtag_break)) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam jtag_break_88.GSR = "ENABLED";
    FD1P3AX jtag_reset_89 (.D(n41399), .SP(w_clk_cpu_enable_271), .CK(w_clk_cpu), 
            .Q(reset_exception)) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam jtag_reset_89.GSR = "ENABLED";
    FD1P3AX uart_rx_byte_i1 (.D(jtag_reg_q[0]), .SP(jrx_csr_read_data_8__N_2865), 
            .CK(w_clk_cpu), .Q(\jrx_csr_read_data[0] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_rx_byte_i1.GSR = "ENABLED";
    FD1S3AX rx_toggle_81 (.D(rx_toggle_N_2930), .CK(jtag_update_N_2932), 
            .Q(rx_toggle)) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(279[4:31])
    defparam rx_toggle_81.GSR = "ENABLED";
    FD1P3AX uart_rx_valid_93 (.D(jrx_csr_read_data_8__N_2865), .SP(w_clk_cpu_enable_275), 
            .CK(w_clk_cpu), .Q(\jtag_reg_addr_d[1] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_rx_valid_93.GSR = "ENABLED";
    FD1P3IX jtag_reg_d_i4 (.D(uart_tx_byte[4]), .SP(w_clk_cpu_enable_872), 
            .CD(GND_net), .CK(w_clk_cpu), .Q(jtag_reg_d[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam jtag_reg_d_i4.GSR = "ENABLED";
    FD1P3IX uart_tx_valid_91 (.D(n42726), .SP(w_clk_cpu_enable_330), .CD(n24867), 
            .CK(w_clk_cpu), .Q(\jtag_reg_addr_d[0] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_tx_valid_91.GSR = "ENABLED";
    FD1P3AX uart_rx_byte_i8 (.D(jtag_reg_q[7]), .SP(jrx_csr_read_data_8__N_2865), 
            .CK(w_clk_cpu), .Q(\jrx_csr_read_data[7] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_rx_byte_i8.GSR = "ENABLED";
    FD1P3AX uart_rx_byte_i7 (.D(jtag_reg_q[6]), .SP(jrx_csr_read_data_8__N_2865), 
            .CK(w_clk_cpu), .Q(\jrx_csr_read_data[6] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_rx_byte_i7.GSR = "ENABLED";
    FD1P3AX uart_rx_byte_i6 (.D(jtag_reg_q[5]), .SP(jrx_csr_read_data_8__N_2865), 
            .CK(w_clk_cpu), .Q(\jrx_csr_read_data[5] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_rx_byte_i6.GSR = "ENABLED";
    FD1P3AX uart_rx_byte_i5 (.D(jtag_reg_q[4]), .SP(jrx_csr_read_data_8__N_2865), 
            .CK(w_clk_cpu), .Q(\jrx_csr_read_data[4] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_rx_byte_i5.GSR = "ENABLED";
    FD1P3AX uart_rx_byte_i4 (.D(jtag_reg_q[3]), .SP(jrx_csr_read_data_8__N_2865), 
            .CK(w_clk_cpu), .Q(\jrx_csr_read_data[3] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_rx_byte_i4.GSR = "ENABLED";
    FD1P3AX uart_rx_byte_i3 (.D(jtag_reg_q[2]), .SP(jrx_csr_read_data_8__N_2865), 
            .CK(w_clk_cpu), .Q(\jrx_csr_read_data[2] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_rx_byte_i3.GSR = "ENABLED";
    FD1P3AX uart_rx_byte_i2 (.D(jtag_reg_q[1]), .SP(jrx_csr_read_data_8__N_2865), 
            .CK(w_clk_cpu), .Q(\jrx_csr_read_data[1] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_rx_byte_i2.GSR = "ENABLED";
    FD1P3IX jtag_reg_d_i0 (.D(uart_tx_byte[0]), .SP(w_clk_cpu_enable_872), 
            .CD(GND_net), .CK(w_clk_cpu), .Q(jtag_reg_d[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam jtag_reg_d_i0.GSR = "ENABLED";
    LUT4 i38031_2_lut_rep_260_3_lut_4_lut_3_lut_3_lut_4_lut (.A(n41428), .B(n39970), 
         .C(cycles_5__N_2495), .Z(w_clk_cpu_enable_865)) /* synthesis lut_function=(!(A (C)+!A !(B+!(C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2421[13:30])
    defparam i38031_2_lut_rep_260_3_lut_4_lut_3_lut_3_lut_4_lut.init = 16'h4f4f;
    LUT4 i38040_2_lut_rep_259_3_lut_4_lut_3_lut_3_lut_4_lut (.A(n41428), .B(n39970), 
         .C(cycles_5__N_2495), .Z(w_clk_cpu_enable_958)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2421[13:30])
    defparam i38040_2_lut_rep_259_3_lut_4_lut_3_lut_3_lut_4_lut.init = 16'h4040;
    LUT4 i37840_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n41428), .B(x_result_sel_csr_d), 
         .C(branch_flushX_m_N_1116), .D(cycles_5__N_2495), .Z(n22501)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2421[13:30])
    defparam i37840_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h4440;
    LUT4 i23501_2_lut_3_lut_4_lut_4_lut_4_lut (.A(n41428), .B(n41417), .C(branch_flushX_m_N_1116), 
         .D(cycles_5__N_2495), .Z(n26142)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2421[13:30])
    defparam i23501_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'h4440;
    LUT4 i37889_2_lut_rep_262_3_lut_4_lut_4_lut_4_lut (.A(n41428), .B(n39970), 
         .C(branch_flushX_m_N_1116), .D(cycles_5__N_2495), .Z(w_clk_cpu_enable_983)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2421[13:30])
    defparam i37889_2_lut_rep_262_3_lut_4_lut_4_lut_4_lut.init = 16'h4440;
    LUT4 n24961_bdd_4_lut_38191 (.A(n41443), .B(jtag_reg_addr_q[1]), .C(jtag_reg_addr_q[2]), 
         .D(jtag_reg_addr_q[0]), .Z(n40543)) /* synthesis lut_function=(!(A (C+(D))+!A ((C+(D))+!B))) */ ;
    defparam n24961_bdd_4_lut_38191.init = 16'h000e;
    LUT4 i3_4_lut (.A(n41484), .B(jtag_reg_q[7]), .C(n41483), .D(n25688), 
         .Z(n38722)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(475[7:15])
    defparam i3_4_lut.init = 16'hffdf;
    LUT4 rx_toggle_I_0_1_lut (.A(rx_toggle), .Z(rx_toggle_N_2930)) /* synthesis lut_function=(!(A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(279[20:30])
    defparam rx_toggle_I_0_1_lut.init = 16'h5555;
    LUT4 i37977_4_lut (.A(\csr_x[0] ), .B(n39169), .C(n38725), .D(n4), 
         .Z(w_clk_cpu_enable_275)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A ((D)+!B))) */ ;
    defparam i37977_4_lut.init = 16'h0ace;
    LUT4 i38024_2_lut_rep_312 (.A(jtag_reg_q[4]), .B(n38722), .Z(n41399)) /* synthesis lut_function=(!((B)+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(424[7] 494[12])
    defparam i38024_2_lut_rep_312.init = 16'h2222;
    LUT4 i1_2_lut_3_lut (.A(jtag_reg_q[4]), .B(n38722), .C(jtag_reg_d_7__N_505), 
         .Z(w_clk_cpu_enable_271)) /* synthesis lut_function=(A ((C)+!B)+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(424[7] 494[12])
    defparam i1_2_lut_3_lut.init = 16'hf2f2;
    LUT4 i38028_2_lut_rep_313 (.A(jtag_reg_q[4]), .B(n38722), .Z(n41400)) /* synthesis lut_function=(!(A+(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(424[7] 494[12])
    defparam i38028_2_lut_rep_313.init = 16'h1111;
    LUT4 i1_2_lut_3_lut_adj_189 (.A(jtag_reg_q[4]), .B(n38722), .C(jtag_reg_d_7__N_505), 
         .Z(w_clk_cpu_enable_270)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(424[7] 494[12])
    defparam i1_2_lut_3_lut_adj_189.init = 16'hf1f1;
    LUT4 i2_4_lut (.A(jtag_reg_addr_q[0]), .B(jtag_reg_addr_q[2]), .C(n10), 
         .D(jtag_reg_addr_q[1]), .Z(w_clk_cpu_enable_872)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2_4_lut.init = 16'h1000;
    LUT4 i24_2_lut (.A(rx_toggle_r_r_r), .B(rx_toggle_r_r), .Z(n10)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i24_2_lut.init = 16'h6666;
    FD1P3AX uart_tx_byte_i0_i7 (.D(\operand_1_x[7] ), .SP(w_clk_cpu_enable_769), 
            .CK(w_clk_cpu), .Q(uart_tx_byte[7])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_tx_byte_i0_i7.GSR = "ENABLED";
    FD1P3AX uart_tx_byte_i0_i6 (.D(\operand_1_x[6] ), .SP(w_clk_cpu_enable_769), 
            .CK(w_clk_cpu), .Q(uart_tx_byte[6])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_tx_byte_i0_i6.GSR = "ENABLED";
    FD1P3AX uart_tx_byte_i0_i5 (.D(\operand_1_x[5] ), .SP(w_clk_cpu_enable_769), 
            .CK(w_clk_cpu), .Q(uart_tx_byte[5])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_tx_byte_i0_i5.GSR = "ENABLED";
    FD1P3AX uart_tx_byte_i0_i4 (.D(\operand_1_x[4] ), .SP(w_clk_cpu_enable_769), 
            .CK(w_clk_cpu), .Q(uart_tx_byte[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_tx_byte_i0_i4.GSR = "ENABLED";
    FD1P3AX uart_tx_byte_i0_i3 (.D(\operand_1_x[3] ), .SP(w_clk_cpu_enable_769), 
            .CK(w_clk_cpu), .Q(uart_tx_byte[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_tx_byte_i0_i3.GSR = "ENABLED";
    FD1P3AX uart_tx_byte_i0_i2 (.D(\operand_1_x[2] ), .SP(w_clk_cpu_enable_769), 
            .CK(w_clk_cpu), .Q(uart_tx_byte[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_tx_byte_i0_i2.GSR = "ENABLED";
    FD1P3AX uart_tx_byte_i0_i1 (.D(\operand_1_x[1] ), .SP(w_clk_cpu_enable_769), 
            .CK(w_clk_cpu), .Q(uart_tx_byte[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam uart_tx_byte_i0_i1.GSR = "ENABLED";
    FD1P3IX jtag_reg_d_i5 (.D(uart_tx_byte[5]), .SP(w_clk_cpu_enable_872), 
            .CD(GND_net), .CK(w_clk_cpu), .Q(jtag_reg_d[5])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=11, LSE_RCOL=6, LSE_LLINE=1163, LSE_RLINE=1208 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(339[4] 584[7])
    defparam jtag_reg_d_i5.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_190 (.A(jtag_reg_addr_q[1]), .B(jtag_reg_addr_q[2]), 
         .C(jtag_reg_addr_q[0]), .Z(n25688)) /* synthesis lut_function=(A+(B+(C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(429[7:15])
    defparam i1_2_lut_3_lut_adj_190.init = 16'hfefe;
    LUT4 i1_3_lut_4_lut (.A(jtag_reg_addr_q[1]), .B(jtag_reg_addr_q[2]), 
         .C(rx_toggle_r_r), .D(rx_toggle_r_r_r), .Z(n4)) /* synthesis lut_function=(A+(B+(C (D)+!C !(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(429[7:15])
    defparam i1_3_lut_4_lut.init = 16'hfeef;
    LUT4 i2_3_lut_4_lut_adj_191 (.A(jtag_reg_addr_q[1]), .B(jtag_reg_addr_q[2]), 
         .C(n41484), .D(jtag_reg_addr_q[0]), .Z(jrx_csr_read_data_8__N_2865)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(429[7:15])
    defparam i2_3_lut_4_lut_adj_191.init = 16'h1000;
    LUT4 i1_2_lut_rep_396 (.A(jtag_reg_q[6]), .B(jtag_reg_q[5]), .Z(n41483)) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(431[5] 466[12])
    defparam i1_2_lut_rep_396.init = 16'h8888;
    LUT4 i36621_2_lut_3_lut_4_lut (.A(jtag_reg_q[6]), .B(jtag_reg_q[5]), 
         .C(jtag_reg_addr_q[0]), .D(jtag_reg_q[7]), .Z(n39169)) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(431[5] 466[12])
    defparam i36621_2_lut_3_lut_4_lut.init = 16'hf0f8;
    LUT4 i2_2_lut_rep_356_3_lut (.A(jtag_reg_q[6]), .B(jtag_reg_q[5]), .C(jtag_reg_q[7]), 
         .Z(n41443)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(431[5] 466[12])
    defparam i2_2_lut_rep_356_3_lut.init = 16'h0808;
    LUT4 rx_toggle_r_r_I_0_2_lut_rep_397 (.A(rx_toggle_r_r), .B(rx_toggle_r_r_r), 
         .Z(n41484)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(424[11:43])
    defparam rx_toggle_r_r_I_0_2_lut_rep_397.init = 16'h6666;
    LUT4 i37974_2_lut_3_lut (.A(rx_toggle_r_r), .B(rx_toggle_r_r_r), .C(n40543), 
         .Z(n24867)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_jtag.v(424[11:43])
    defparam i37974_2_lut_3_lut.init = 16'h6060;
    
endmodule
//
// Verilog Description of module lm32_interrupt
//

module lm32_interrupt (im, w_clk_cpu, operand_1_x, \im[18] , \im[17] , 
            \im[16] , \im[15] , \im[14] , \im[13] , \im[12] , \im[11] , 
            \im[10] , \im[9] , \im[31] , \im[8] , \im[30] , \im[7] , 
            \im[29] , \im[6] , \im[28] , \im[5] , bie, bie_N_2835, 
            \im[27] , \im[4] , eie, n23750, ie, \csr_x[0] , n21263, 
            \im[26] , \im[3] , n41474, \csr_x[1] , n25705, \im[25] , 
            \im[2] , \im[24] , \im[1] , \im[23] , n41473, n41472, 
            n25625, bret_q_x, w_clk_cpu_enable_984, n4, jtag_reg_d_7__N_505, 
            n41359, ie_N_2822, n41357, n41502, \csr_x[2] , n38725, 
            \im[22] , w_clk_cpu_enable_330, n41391, eret_x, bret_x, 
            n41351, ie_N_2821) /* synthesis syn_module_defined=1 */ ;
    output [31:0]im;
    input w_clk_cpu;
    input [31:0]operand_1_x;
    output \im[18] ;
    output \im[17] ;
    output \im[16] ;
    output \im[15] ;
    output \im[14] ;
    output \im[13] ;
    output \im[12] ;
    output \im[11] ;
    output \im[10] ;
    output \im[9] ;
    output \im[31] ;
    output \im[8] ;
    output \im[30] ;
    output \im[7] ;
    output \im[29] ;
    output \im[6] ;
    output \im[28] ;
    output \im[5] ;
    output bie;
    input bie_N_2835;
    output \im[27] ;
    output \im[4] ;
    output eie;
    input n23750;
    output ie;
    input \csr_x[0] ;
    output n21263;
    output \im[26] ;
    output \im[3] ;
    input n41474;
    input \csr_x[1] ;
    output n25705;
    output \im[25] ;
    output \im[2] ;
    output \im[24] ;
    output \im[1] ;
    output \im[23] ;
    input n41473;
    input n41472;
    output n25625;
    input bret_q_x;
    input w_clk_cpu_enable_984;
    input n4;
    input jtag_reg_d_7__N_505;
    input n41359;
    output ie_N_2822;
    input n41357;
    input n41502;
    input \csr_x[2] ;
    output n38725;
    output \im[22] ;
    output w_clk_cpu_enable_330;
    input n41391;
    input eret_x;
    input bret_x;
    input n41351;
    input ie_N_2821;
    
    wire w_clk_cpu /* synthesis SET_AS_NETWORK=w_clk_cpu, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(22[6:15])
    
    wire w_clk_cpu_enable_709;
    wire [31:0]im_c;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(141[22:24])
    
    wire w_clk_cpu_enable_255, w_clk_cpu_enable_273, w_clk_cpu_enable_982, 
        n4_adj_3698;
    
    FD1P3AX im_i0_i21 (.D(operand_1_x[21]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(im[21])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i21.GSR = "ENABLED";
    FD1P3AX im_i0_i20 (.D(operand_1_x[20]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(im[20])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i20.GSR = "ENABLED";
    FD1P3AX im_i0_i19 (.D(operand_1_x[19]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(im[19])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i19.GSR = "ENABLED";
    FD1P3AX im_i0_i0 (.D(operand_1_x[0]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(im_c[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i0.GSR = "ENABLED";
    FD1P3AX im_i0_i18 (.D(operand_1_x[18]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[18] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i18.GSR = "ENABLED";
    FD1P3AX im_i0_i17 (.D(operand_1_x[17]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[17] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i17.GSR = "ENABLED";
    FD1P3AX im_i0_i16 (.D(operand_1_x[16]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[16] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i16.GSR = "ENABLED";
    FD1P3AX im_i0_i15 (.D(operand_1_x[15]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[15] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i15.GSR = "ENABLED";
    FD1P3AX im_i0_i14 (.D(operand_1_x[14]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[14] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i14.GSR = "ENABLED";
    FD1P3AX im_i0_i13 (.D(operand_1_x[13]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[13] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i13.GSR = "ENABLED";
    FD1P3AX im_i0_i12 (.D(operand_1_x[12]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[12] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i12.GSR = "ENABLED";
    FD1P3AX im_i0_i11 (.D(operand_1_x[11]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[11] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i11.GSR = "ENABLED";
    FD1P3AX im_i0_i10 (.D(operand_1_x[10]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[10] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i10.GSR = "ENABLED";
    FD1P3AX im_i0_i9 (.D(operand_1_x[9]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[9] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i9.GSR = "ENABLED";
    FD1P3AX im_i0_i31 (.D(operand_1_x[31]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[31] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i31.GSR = "ENABLED";
    FD1P3AX im_i0_i8 (.D(operand_1_x[8]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[8] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i8.GSR = "ENABLED";
    FD1P3AX im_i0_i30 (.D(operand_1_x[30]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[30] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i30.GSR = "ENABLED";
    FD1P3AX im_i0_i7 (.D(operand_1_x[7]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[7] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i7.GSR = "ENABLED";
    FD1P3AX im_i0_i29 (.D(operand_1_x[29]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[29] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i29.GSR = "ENABLED";
    FD1P3AX im_i0_i6 (.D(operand_1_x[6]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[6] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i6.GSR = "ENABLED";
    FD1P3AX im_i0_i28 (.D(operand_1_x[28]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[28] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i28.GSR = "ENABLED";
    FD1P3AX im_i0_i5 (.D(operand_1_x[5]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[5] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i5.GSR = "ENABLED";
    FD1P3AX bie_68 (.D(bie_N_2835), .SP(w_clk_cpu_enable_255), .CK(w_clk_cpu), 
            .Q(bie));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam bie_68.GSR = "ENABLED";
    FD1P3AX im_i0_i27 (.D(operand_1_x[27]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[27] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i27.GSR = "ENABLED";
    FD1P3AX im_i0_i4 (.D(operand_1_x[4]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[4] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i4.GSR = "ENABLED";
    FD1P3AX eie_67 (.D(n23750), .SP(w_clk_cpu_enable_273), .CK(w_clk_cpu), 
            .Q(eie));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam eie_67.GSR = "ENABLED";
    LUT4 mux_19115_Mux_0_i1_3_lut (.A(ie), .B(im_c[0]), .C(\csr_x[0] ), 
         .Z(n21263)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(173[5] 186[12])
    defparam mux_19115_Mux_0_i1_3_lut.init = 16'hcaca;
    FD1P3AX im_i0_i26 (.D(operand_1_x[26]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[26] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i26.GSR = "ENABLED";
    FD1P3AX im_i0_i3 (.D(operand_1_x[3]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[3] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i3.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut (.A(\csr_x[0] ), .B(n41474), .C(\csr_x[1] ), .Z(n25705)) /* synthesis lut_function=(A+(B+(C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(183[5:17])
    defparam i1_2_lut_3_lut.init = 16'hfefe;
    FD1P3AX im_i0_i25 (.D(operand_1_x[25]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[25] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i25.GSR = "ENABLED";
    FD1P3AX im_i0_i2 (.D(operand_1_x[2]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[2] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i2.GSR = "ENABLED";
    FD1P3AX im_i0_i24 (.D(operand_1_x[24]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[24] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i24.GSR = "ENABLED";
    FD1P3AX im_i0_i1 (.D(operand_1_x[1]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[1] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i1.GSR = "ENABLED";
    FD1P3AX im_i0_i23 (.D(operand_1_x[23]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[23] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i23.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(n25705), .B(n41473), .C(n41472), .D(n25625), .Z(w_clk_cpu_enable_255)) /* synthesis lut_function=(!(A (B+!(C))+!A (B+!(C+(D))))) */ ;
    defparam i1_4_lut.init = 16'h3130;
    LUT4 i29899_4_lut (.A(bret_q_x), .B(w_clk_cpu_enable_984), .C(n4), 
         .D(jtag_reg_d_7__N_505), .Z(w_clk_cpu_enable_982)) /* synthesis lut_function=(A (B+(D))+!A (B (C)+!B (C (D)))) */ ;
    defparam i29899_4_lut.init = 16'hfac8;
    LUT4 ie_I_111_4_lut (.A(operand_1_x[0]), .B(bie), .C(bret_q_x), .D(n41359), 
         .Z(ie_N_2822)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(266[18] 281[16])
    defparam ie_I_111_4_lut.init = 16'hcac0;
    LUT4 i2_4_lut (.A(\csr_x[1] ), .B(n41357), .C(n41502), .D(\csr_x[2] ), 
         .Z(n38725)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(183[5:17])
    defparam i2_4_lut.init = 16'hf7ff;
    LUT4 i1_3_lut_4_lut (.A(n25625), .B(n41472), .C(n41473), .D(n25705), 
         .Z(w_clk_cpu_enable_273)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(242[14] 282[12])
    defparam i1_3_lut_4_lut.init = 16'hf0f2;
    FD1P3AX im_i0_i22 (.D(operand_1_x[22]), .SP(w_clk_cpu_enable_709), .CK(w_clk_cpu), 
            .Q(\im[22] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=1133, LSE_RLINE=1158 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam im_i0_i22.GSR = "ENABLED";
    LUT4 i38017_2_lut (.A(\csr_x[0] ), .B(n38725), .Z(w_clk_cpu_enable_330)) /* synthesis lut_function=(!(A+(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(183[5:17])
    defparam i38017_2_lut.init = 16'h1111;
    LUT4 i2_4_lut_adj_186 (.A(n41357), .B(n41391), .C(eret_x), .D(bret_x), 
         .Z(n25625)) /* synthesis lut_function=(!((B (C+(D)))+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(242[14] 282[12])
    defparam i2_4_lut_adj_186.init = 16'h222a;
    LUT4 i1_4_lut_adj_187 (.A(n41474), .B(n41351), .C(n41473), .D(n4_adj_3698), 
         .Z(w_clk_cpu_enable_709)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(242[14] 282[12])
    defparam i1_4_lut_adj_187.init = 16'h0004;
    LUT4 i1_2_lut (.A(\csr_x[1] ), .B(\csr_x[0] ), .Z(n4_adj_3698)) /* synthesis lut_function=(A+!(B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(184[5:17])
    defparam i1_2_lut.init = 16'hbbbb;
    FD1P3IX ie_66 (.D(ie_N_2821), .SP(w_clk_cpu_enable_982), .CD(jtag_reg_d_7__N_505), 
            .CK(w_clk_cpu), .Q(ie));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_interrupt.v(232[5] 283[8])
    defparam ie_66.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module lm32_instruction_unit
//

module lm32_instruction_unit (pc_d, w_clk_cpu, w_clk_cpu_enable_983, pc_f, 
            \instruction_d[13] , w_clk_cpu_enable_984, branch_taken_m, 
            w_clk_cpu_enable_914, \instruction_d[12] , \instruction_d[11] , 
            \instruction_d[10] , \instruction_d[9] , \instruction_d[8] , 
            \instruction_d[7] , \instruction_d[6] , \instruction_d[5] , 
            \instruction_d[4] , \instruction_d[3] , \instruction_d[2] , 
            GND_net, pc_m, w_clk_cpu_enable_972, \LM32I_ADR_O[2] , w_clk_cpu_enable_763, 
            SHAREDBUS_DAT_O, LM32I_CYC_O, n37179, \instruction_d[0] , 
            \selected_1__N_344[0] , w_clk_cpu_enable_216, \instruction_d[1] , 
            n41375, n41504, \branch_target_d[3] , n42746, n41459, 
            branch_target_m, i_cyc_o_N_1759, valid_d, n41394, \LM32I_ADR_O[31] , 
            bus_error_f_N_1764, \LM32I_ADR_O[30] , \branch_target_d[30] , 
            \branch_target_d[31] , \LM32I_ADR_O[29] , \branch_target_d[28] , 
            \branch_target_d[29] , \LM32I_ADR_O[28] , \branch_target_d[26] , 
            \branch_target_d[27] , \LM32I_ADR_O[27] , \branch_target_d[24] , 
            \branch_target_d[25] , \LM32I_ADR_O[26] , \LM32I_ADR_O[25] , 
            \branch_target_d[22] , \branch_target_d[23] , \branch_target_d[20] , 
            \branch_target_d[21] , \LM32I_ADR_O[24] , \LM32I_ADR_O[23] , 
            \branch_target_d[18] , \branch_target_d[19] , \branch_target_d[16] , 
            \branch_target_d[17] , \LM32I_ADR_O[22] , \branch_target_d[14] , 
            \branch_target_d[15] , \LM32I_ADR_O[21] , \branch_target_d[12] , 
            \branch_target_d[13] , \LM32I_ADR_O[20] , \LM32I_ADR_O[19] , 
            \LM32I_ADR_O[18] , \LM32I_ADR_O[17] , \branch_target_d[6] , 
            \branch_target_d[7] , \LM32I_ADR_O[16] , \LM32I_ADR_O[15] , 
            \LM32I_ADR_O[14] , \branch_target_d[8] , \branch_target_d[9] , 
            \LM32I_ADR_O[13] , \LM32I_ADR_O[12] , \branch_target_d[4] , 
            \branch_target_d[5] , \LM32I_ADR_O[11] , \branch_target_d[10] , 
            \branch_target_d[11] , \LM32I_ADR_O[10] , \LM32I_ADR_O[9] , 
            \LM32I_ADR_O[8] , \LM32I_ADR_O[7] , \LM32I_ADR_O[6] , \LM32I_ADR_O[5] , 
            \LM32I_ADR_O[4] , \LM32I_ADR_O[3] , n42740, n41479, n38871, 
            w_clk_cpu_enable_878, bus_error_d, \instruction_d[31] , \instruction_d[30] , 
            \logic_op_d[3] , sign_extend_d, size_d, read_idx_0_d, w_clk_cpu_enable_985, 
            read_idx_1_d, \instruction_d[15] , \instruction_d[14] ) /* synthesis syn_module_defined=1 */ ;
    output [31:2]pc_d;
    input w_clk_cpu;
    input w_clk_cpu_enable_983;
    output [31:2]pc_f;
    output \instruction_d[13] ;
    input w_clk_cpu_enable_984;
    input branch_taken_m;
    input w_clk_cpu_enable_914;
    output \instruction_d[12] ;
    output \instruction_d[11] ;
    output \instruction_d[10] ;
    output \instruction_d[9] ;
    output \instruction_d[8] ;
    output \instruction_d[7] ;
    output \instruction_d[6] ;
    output \instruction_d[5] ;
    output \instruction_d[4] ;
    output \instruction_d[3] ;
    output \instruction_d[2] ;
    input GND_net;
    output [31:2]pc_m;
    input w_clk_cpu_enable_972;
    output \LM32I_ADR_O[2] ;
    input w_clk_cpu_enable_763;
    input [31:0]SHAREDBUS_DAT_O;
    output LM32I_CYC_O;
    input n37179;
    output \instruction_d[0] ;
    output \selected_1__N_344[0] ;
    input w_clk_cpu_enable_216;
    output \instruction_d[1] ;
    input n41375;
    input n41504;
    input \branch_target_d[3] ;
    input n42746;
    input n41459;
    input [31:2]branch_target_m;
    input i_cyc_o_N_1759;
    input valid_d;
    input n41394;
    output \LM32I_ADR_O[31] ;
    input bus_error_f_N_1764;
    output \LM32I_ADR_O[30] ;
    input \branch_target_d[30] ;
    input \branch_target_d[31] ;
    output \LM32I_ADR_O[29] ;
    input \branch_target_d[28] ;
    input \branch_target_d[29] ;
    output \LM32I_ADR_O[28] ;
    input \branch_target_d[26] ;
    input \branch_target_d[27] ;
    output \LM32I_ADR_O[27] ;
    input \branch_target_d[24] ;
    input \branch_target_d[25] ;
    output \LM32I_ADR_O[26] ;
    output \LM32I_ADR_O[25] ;
    input \branch_target_d[22] ;
    input \branch_target_d[23] ;
    input \branch_target_d[20] ;
    input \branch_target_d[21] ;
    output \LM32I_ADR_O[24] ;
    output \LM32I_ADR_O[23] ;
    input \branch_target_d[18] ;
    input \branch_target_d[19] ;
    input \branch_target_d[16] ;
    input \branch_target_d[17] ;
    output \LM32I_ADR_O[22] ;
    input \branch_target_d[14] ;
    input \branch_target_d[15] ;
    output \LM32I_ADR_O[21] ;
    input \branch_target_d[12] ;
    input \branch_target_d[13] ;
    output \LM32I_ADR_O[20] ;
    output \LM32I_ADR_O[19] ;
    output \LM32I_ADR_O[18] ;
    output \LM32I_ADR_O[17] ;
    input \branch_target_d[6] ;
    input \branch_target_d[7] ;
    output \LM32I_ADR_O[16] ;
    output \LM32I_ADR_O[15] ;
    output \LM32I_ADR_O[14] ;
    input \branch_target_d[8] ;
    input \branch_target_d[9] ;
    output \LM32I_ADR_O[13] ;
    output \LM32I_ADR_O[12] ;
    input \branch_target_d[4] ;
    input \branch_target_d[5] ;
    output \LM32I_ADR_O[11] ;
    input \branch_target_d[10] ;
    input \branch_target_d[11] ;
    output \LM32I_ADR_O[10] ;
    output \LM32I_ADR_O[9] ;
    output \LM32I_ADR_O[8] ;
    output \LM32I_ADR_O[7] ;
    output \LM32I_ADR_O[6] ;
    output \LM32I_ADR_O[5] ;
    output \LM32I_ADR_O[4] ;
    output \LM32I_ADR_O[3] ;
    input n42740;
    input n41479;
    input n38871;
    input w_clk_cpu_enable_878;
    output bus_error_d;
    output \instruction_d[31] ;
    output \instruction_d[30] ;
    output \logic_op_d[3] ;
    output sign_extend_d;
    output [1:0]size_d;
    output [4:0]read_idx_0_d;
    input w_clk_cpu_enable_985;
    output [4:0]read_idx_1_d;
    output \instruction_d[15] ;
    output \instruction_d[14] ;
    
    wire w_clk_cpu /* synthesis SET_AS_NETWORK=w_clk_cpu, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(22[6:15])
    wire [31:0]wb_data_f;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(352[29:38])
    wire [31:2]pc_x;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(633[21:25])
    wire [29:0]pc_a_31__N_1556;
    wire [29:0]pc_a_31__N_1586;
    wire [31:2]pc_a;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(334[20:24])
    
    wire n36607, n22255, n22254, n36608, w_clk_cpu_enable_558, i_cyc_o_N_1754, 
        n36606, n22257, n22256, n36583, n22272, n22271, n36584, 
        n36605, n22259, n22258, n36604, n22261, n22260, n36603, 
        n22263, n22262, n36602, n22265, n22264, n36601, n22267, 
        n22266, n36600, n22269, n22268, n36599, n22270, bus_error_f, 
        w_clk_cpu_enable_587, n36597, n22244, n22243, n36596, n22246, 
        n22245, n36595, n22248, n22247, n36594, n22250, n22249, 
        n36593, n22252, n22251, n36592, n22253, n36591, n36590, 
        n36589, n36588, n36585, n36586, n36613, n36612, n36611, 
        n36610, n36609, n36587;
    
    FD1P3AX pc_d_i2_i14 (.D(pc_f[14]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_d[14])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i14.GSR = "ENABLED";
    FD1P3AX pc_d_i2_i13 (.D(pc_f[13]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_d[13])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i13.GSR = "ENABLED";
    FD1P3AX pc_d_i2_i31 (.D(pc_f[31]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_d[31])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i31.GSR = "ENABLED";
    FD1P3AX pc_d_i2_i12 (.D(pc_f[12]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_d[12])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i12.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i13 (.D(wb_data_f[13]), .SP(w_clk_cpu_enable_983), 
            .CK(w_clk_cpu), .Q(\instruction_d[13] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i13.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i17 (.D(pc_d[17]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[17])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i17.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i16 (.D(pc_d[16]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[16])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i16.GSR = "ENABLED";
    FD1P3AX pc_d_i2_i2 (.D(pc_f[2]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_d[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i2.GSR = "ENABLED";
    FD1P3AX pc_d_i2_i30 (.D(pc_f[30]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_d[30])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i30.GSR = "ENABLED";
    FD1P3AX pc_d_i2_i11 (.D(pc_f[11]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_d[11])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i11.GSR = "ENABLED";
    FD1P3AX pc_d_i2_i29 (.D(pc_f[29]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_d[29])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i29.GSR = "ENABLED";
    LUT4 pc_a_31__I_0_i29_3_lut (.A(pc_a_31__N_1556[28]), .B(pc_a_31__N_1586[28]), 
         .C(branch_taken_m), .Z(pc_a[30])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i29_3_lut.init = 16'hcaca;
    FD1P3AX pc_d_i2_i28 (.D(pc_f[28]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_d[28])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i28.GSR = "ENABLED";
    FD1P3AX pc_d_i2_i10 (.D(pc_f[10]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_d[10])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i10.GSR = "ENABLED";
    FD1P3AX pc_d_i2_i27 (.D(pc_f[27]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_d[27])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i27.GSR = "ENABLED";
    FD1P3AX pc_d_i2_i9 (.D(pc_f[9]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_d[9])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i9.GSR = "ENABLED";
    FD1P3AX pc_d_i2_i8 (.D(pc_f[8]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_d[8])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i8.GSR = "ENABLED";
    FD1P3AX pc_d_i2_i26 (.D(pc_f[26]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_d[26])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i26.GSR = "ENABLED";
    FD1P3AX pc_d_i2_i7 (.D(pc_f[7]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_d[7])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i7.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i12 (.D(wb_data_f[12]), .SP(w_clk_cpu_enable_914), 
            .CK(w_clk_cpu), .Q(\instruction_d[12] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i12.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i15 (.D(pc_d[15]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[15])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i15.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i14 (.D(pc_d[14]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[14])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i14.GSR = "ENABLED";
    LUT4 pc_a_31__I_0_i28_3_lut (.A(pc_a_31__N_1556[27]), .B(pc_a_31__N_1586[27]), 
         .C(branch_taken_m), .Z(pc_a[29])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i28_3_lut.init = 16'hcaca;
    FD1P3AX instruction_d_i0_i11 (.D(wb_data_f[11]), .SP(w_clk_cpu_enable_914), 
            .CK(w_clk_cpu), .Q(\instruction_d[11] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i11.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i13 (.D(pc_d[13]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[13])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i13.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i12 (.D(pc_d[12]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[12])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i12.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i10 (.D(wb_data_f[10]), .SP(w_clk_cpu_enable_914), 
            .CK(w_clk_cpu), .Q(\instruction_d[10] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i10.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i11 (.D(pc_d[11]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[11])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i11.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i10 (.D(pc_d[10]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[10])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i10.GSR = "ENABLED";
    FD1P3AX pc_d_i2_i6 (.D(pc_f[6]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_d[6])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i6.GSR = "ENABLED";
    LUT4 pc_a_31__I_0_i27_3_lut (.A(pc_a_31__N_1556[26]), .B(pc_a_31__N_1586[26]), 
         .C(branch_taken_m), .Z(pc_a[28])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i27_3_lut.init = 16'hcaca;
    FD1P3AX instruction_d_i0_i9 (.D(wb_data_f[9]), .SP(w_clk_cpu_enable_914), 
            .CK(w_clk_cpu), .Q(\instruction_d[9] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i9.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i9 (.D(pc_d[9]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[9])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i9.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i8 (.D(pc_d[8]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[8])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i8.GSR = "ENABLED";
    LUT4 pc_a_31__I_0_i26_3_lut (.A(pc_a_31__N_1556[25]), .B(pc_a_31__N_1586[25]), 
         .C(branch_taken_m), .Z(pc_a[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i26_3_lut.init = 16'hcaca;
    FD1P3AX instruction_d_i0_i8 (.D(wb_data_f[8]), .SP(w_clk_cpu_enable_914), 
            .CK(w_clk_cpu), .Q(\instruction_d[8] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i8.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i7 (.D(pc_d[7]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[7])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i7.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i6 (.D(pc_d[6]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[6])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i6.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i7 (.D(wb_data_f[7]), .SP(w_clk_cpu_enable_914), 
            .CK(w_clk_cpu), .Q(\instruction_d[7] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i7.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i5 (.D(pc_d[5]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[5])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i5.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i4 (.D(pc_d[4]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i4.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i6 (.D(wb_data_f[6]), .SP(w_clk_cpu_enable_914), 
            .CK(w_clk_cpu), .Q(\instruction_d[6] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i6.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i3 (.D(pc_d[3]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i3.GSR = "ENABLED";
    LUT4 pc_a_31__I_0_i25_3_lut (.A(pc_a_31__N_1556[24]), .B(pc_a_31__N_1586[24]), 
         .C(branch_taken_m), .Z(pc_a[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i25_3_lut.init = 16'hcaca;
    FD1P3AX instruction_d_i0_i5 (.D(wb_data_f[5]), .SP(w_clk_cpu_enable_914), 
            .CK(w_clk_cpu), .Q(\instruction_d[5] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i5.GSR = "ENABLED";
    LUT4 pc_a_31__I_0_i24_3_lut (.A(pc_a_31__N_1556[23]), .B(pc_a_31__N_1586[23]), 
         .C(branch_taken_m), .Z(pc_a[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i24_3_lut.init = 16'hcaca;
    FD1P3AX instruction_d_i0_i4 (.D(wb_data_f[4]), .SP(w_clk_cpu_enable_983), 
            .CK(w_clk_cpu), .Q(\instruction_d[4] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i4.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i3 (.D(wb_data_f[3]), .SP(w_clk_cpu_enable_983), 
            .CK(w_clk_cpu), .Q(\instruction_d[3] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i3.GSR = "ENABLED";
    FD1P3AX pc_d_i2_i25 (.D(pc_f[25]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_d[25])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i25.GSR = "ENABLED";
    LUT4 pc_a_31__I_0_i23_3_lut (.A(pc_a_31__N_1556[22]), .B(pc_a_31__N_1586[22]), 
         .C(branch_taken_m), .Z(pc_a[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i23_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_0_i22_3_lut (.A(pc_a_31__N_1556[21]), .B(pc_a_31__N_1586[21]), 
         .C(branch_taken_m), .Z(pc_a[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i22_3_lut.init = 16'hcaca;
    FD1P3AX instruction_d_i0_i2 (.D(wb_data_f[2]), .SP(w_clk_cpu_enable_983), 
            .CK(w_clk_cpu), .Q(\instruction_d[2] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i2.GSR = "ENABLED";
    FD1P3AX pc_d_i2_i5 (.D(pc_f[5]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_d[5])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i5.GSR = "ENABLED";
    CCU2D add_18875_rep_2_19 (.A0(pc_f[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pc_f[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n36607), .COUT(n36608), .S0(n22255), .S1(n22254));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_2_19.INIT0 = 16'hfaaa;
    defparam add_18875_rep_2_19.INIT1 = 16'hfaaa;
    defparam add_18875_rep_2_19.INJECT1_0 = "NO";
    defparam add_18875_rep_2_19.INJECT1_1 = "NO";
    LUT4 pc_a_31__I_0_i21_3_lut (.A(pc_a_31__N_1556[20]), .B(pc_a_31__N_1586[20]), 
         .C(branch_taken_m), .Z(pc_a[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i21_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_0_i20_3_lut (.A(pc_a_31__N_1556[19]), .B(pc_a_31__N_1586[19]), 
         .C(branch_taken_m), .Z(pc_a[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i20_3_lut.init = 16'hcaca;
    FD1P3AX pc_d_i2_i24 (.D(pc_f[24]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_d[24])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i24.GSR = "ENABLED";
    FD1P3AX pc_d_i2_i4 (.D(pc_f[4]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_d[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i4.GSR = "ENABLED";
    LUT4 pc_a_31__I_0_i19_3_lut (.A(pc_a_31__N_1556[18]), .B(pc_a_31__N_1586[18]), 
         .C(branch_taken_m), .Z(pc_a[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i19_3_lut.init = 16'hcaca;
    FD1P3AX pc_d_i2_i23 (.D(pc_f[23]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_d[23])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i23.GSR = "ENABLED";
    FD1P3AX pc_d_i2_i3 (.D(pc_f[3]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_d[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i3.GSR = "ENABLED";
    LUT4 pc_a_31__I_0_i18_3_lut (.A(pc_a_31__N_1556[17]), .B(pc_a_31__N_1586[17]), 
         .C(branch_taken_m), .Z(pc_a[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i18_3_lut.init = 16'hcaca;
    FD1P3AX pc_d_i2_i22 (.D(pc_f[22]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_d[22])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i22.GSR = "ENABLED";
    LUT4 pc_a_31__I_0_i17_3_lut (.A(pc_a_31__N_1556[16]), .B(pc_a_31__N_1586[16]), 
         .C(branch_taken_m), .Z(pc_a[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i17_3_lut.init = 16'hcaca;
    FD1P3AX pc_x_i2_i2 (.D(pc_d[2]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i2.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i2 (.D(pc_x[2]), .SP(w_clk_cpu_enable_972), .CK(w_clk_cpu), 
            .Q(pc_m[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i2.GSR = "ENABLED";
    FD1P3AX i_adr_o__i1 (.D(pc_a[2]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[2] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i1.GSR = "ENABLED";
    FD1P3AX wb_data_f_i0_i0 (.D(SHAREDBUS_DAT_O[0]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i0.GSR = "ENABLED";
    FD1S3AX i_cyc_o_70 (.D(n37179), .CK(w_clk_cpu), .Q(LM32I_CYC_O)) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_cyc_o_70.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i0 (.D(wb_data_f[0]), .SP(w_clk_cpu_enable_983), 
            .CK(w_clk_cpu), .Q(\instruction_d[0] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i0.GSR = "ENABLED";
    FD1P3AX i_stb_o_71 (.D(i_cyc_o_N_1754), .SP(w_clk_cpu_enable_216), .CK(w_clk_cpu), 
            .Q(\selected_1__N_344[0] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_stb_o_71.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i2 (.D(pc_a[2]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_f[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i2.GSR = "ENABLED";
    FD1P3AX pc_d_i2_i21 (.D(pc_f[21]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_d[21])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i21.GSR = "ENABLED";
    FD1P3AX pc_d_i2_i20 (.D(pc_f[20]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_d[20])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i20.GSR = "ENABLED";
    CCU2D add_18875_rep_2_17 (.A0(pc_f[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pc_f[18]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n36606), .COUT(n36607), .S0(n22257), .S1(n22256));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_2_17.INIT0 = 16'hfaaa;
    defparam add_18875_rep_2_17.INIT1 = 16'hfaaa;
    defparam add_18875_rep_2_17.INJECT1_0 = "NO";
    defparam add_18875_rep_2_17.INJECT1_1 = "NO";
    LUT4 pc_a_31__I_0_i16_3_lut (.A(pc_a_31__N_1556[15]), .B(pc_a_31__N_1586[15]), 
         .C(branch_taken_m), .Z(pc_a[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i16_3_lut.init = 16'hcaca;
    FD1P3AX pc_d_i2_i19 (.D(pc_f[19]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_d[19])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i19.GSR = "ENABLED";
    LUT4 pc_a_31__I_0_i15_3_lut (.A(pc_a_31__N_1556[14]), .B(pc_a_31__N_1586[14]), 
         .C(branch_taken_m), .Z(pc_a[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i15_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_0_i14_3_lut (.A(pc_a_31__N_1556[13]), .B(pc_a_31__N_1586[13]), 
         .C(branch_taken_m), .Z(pc_a[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i14_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_0_i13_3_lut (.A(pc_a_31__N_1556[12]), .B(pc_a_31__N_1586[12]), 
         .C(branch_taken_m), .Z(pc_a[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i13_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_0_i12_3_lut (.A(pc_a_31__N_1556[11]), .B(pc_a_31__N_1586[11]), 
         .C(branch_taken_m), .Z(pc_a[13])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i12_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_0_i11_3_lut (.A(pc_a_31__N_1556[10]), .B(pc_a_31__N_1586[10]), 
         .C(branch_taken_m), .Z(pc_a[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i11_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_0_i10_3_lut (.A(pc_a_31__N_1556[9]), .B(pc_a_31__N_1586[9]), 
         .C(branch_taken_m), .Z(pc_a[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i10_3_lut.init = 16'hcaca;
    FD1P3AX instruction_d_i0_i1 (.D(wb_data_f[1]), .SP(w_clk_cpu_enable_914), 
            .CK(w_clk_cpu), .Q(\instruction_d[1] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i1.GSR = "ENABLED";
    LUT4 pc_a_31__I_0_i9_3_lut (.A(pc_a_31__N_1556[8]), .B(pc_a_31__N_1586[8]), 
         .C(branch_taken_m), .Z(pc_a[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i9_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_0_i8_3_lut (.A(pc_a_31__N_1556[7]), .B(pc_a_31__N_1586[7]), 
         .C(branch_taken_m), .Z(pc_a[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i8_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_0_i7_3_lut (.A(pc_a_31__N_1556[6]), .B(pc_a_31__N_1586[6]), 
         .C(branch_taken_m), .Z(pc_a[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i7_3_lut.init = 16'hcaca;
    FD1P3AX pc_d_i2_i18 (.D(pc_f[18]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_d[18])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i18.GSR = "ENABLED";
    LUT4 pc_a_31__I_0_i6_3_lut (.A(pc_a_31__N_1556[5]), .B(pc_a_31__N_1586[5]), 
         .C(branch_taken_m), .Z(pc_a[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i6_3_lut.init = 16'hcaca;
    FD1P3AX pc_d_i2_i17 (.D(pc_f[17]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_d[17])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i17.GSR = "ENABLED";
    LUT4 pc_a_31__I_0_i5_3_lut (.A(pc_a_31__N_1556[4]), .B(pc_a_31__N_1586[4]), 
         .C(branch_taken_m), .Z(pc_a[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i5_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_0_i4_3_lut (.A(pc_a_31__N_1556[3]), .B(pc_a_31__N_1586[3]), 
         .C(branch_taken_m), .Z(pc_a[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i4_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_0_i3_3_lut (.A(pc_a_31__N_1556[2]), .B(pc_a_31__N_1586[2]), 
         .C(branch_taken_m), .Z(pc_a[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i3_3_lut.init = 16'hcaca;
    LUT4 pc_a_31__I_0_i2_3_lut (.A(pc_a_31__N_1556[1]), .B(pc_a_31__N_1586[1]), 
         .C(branch_taken_m), .Z(pc_a[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i2_3_lut.init = 16'hcaca;
    FD1P3AX wb_data_f_i0_i31 (.D(SHAREDBUS_DAT_O[31]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[31])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i31.GSR = "ENABLED";
    FD1P3AX wb_data_f_i0_i30 (.D(SHAREDBUS_DAT_O[30]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[30])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i30.GSR = "ENABLED";
    FD1P3AX wb_data_f_i0_i29 (.D(SHAREDBUS_DAT_O[29]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[29])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i29.GSR = "ENABLED";
    FD1P3AX wb_data_f_i0_i28 (.D(SHAREDBUS_DAT_O[28]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[28])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i28.GSR = "ENABLED";
    FD1P3AX wb_data_f_i0_i27 (.D(SHAREDBUS_DAT_O[27]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[27])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i27.GSR = "ENABLED";
    FD1P3AX wb_data_f_i0_i26 (.D(SHAREDBUS_DAT_O[26]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[26])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i26.GSR = "ENABLED";
    FD1P3AX wb_data_f_i0_i25 (.D(SHAREDBUS_DAT_O[25]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[25])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i25.GSR = "ENABLED";
    FD1P3AX wb_data_f_i0_i24 (.D(SHAREDBUS_DAT_O[24]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[24])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i24.GSR = "ENABLED";
    FD1P3AX wb_data_f_i0_i23 (.D(SHAREDBUS_DAT_O[23]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[23])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i23.GSR = "ENABLED";
    CCU2D add_18875_rep_3_3 (.A0(n22272), .B0(n41375), .C0(n41504), .D0(GND_net), 
          .A1(n22271), .B1(n41375), .C1(\branch_target_d[3] ), .D1(GND_net), 
          .CIN(n36583), .COUT(n36584), .S0(pc_a_31__N_1556[0]), .S1(pc_a_31__N_1556[1]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_3_3.INIT0 = 16'hd2e2;
    defparam add_18875_rep_3_3.INIT1 = 16'hd2e2;
    defparam add_18875_rep_3_3.INJECT1_0 = "NO";
    defparam add_18875_rep_3_3.INJECT1_1 = "NO";
    FD1P3AX wb_data_f_i0_i22 (.D(SHAREDBUS_DAT_O[22]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[22])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i22.GSR = "ENABLED";
    FD1P3AX wb_data_f_i0_i21 (.D(SHAREDBUS_DAT_O[21]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[21])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i21.GSR = "ENABLED";
    LUT4 branch_target_m_31__I_0_i1_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[2]), .D(branch_target_m[2]), .Z(pc_a_31__N_1586[0])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i1_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i30_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[31]), .D(branch_target_m[31]), .Z(pc_a_31__N_1586[29])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i30_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i29_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[30]), .D(branch_target_m[30]), .Z(pc_a_31__N_1586[28])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i29_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i28_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[29]), .D(branch_target_m[29]), .Z(pc_a_31__N_1586[27])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i28_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i27_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[28]), .D(branch_target_m[28]), .Z(pc_a_31__N_1586[26])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i27_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i26_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[27]), .D(branch_target_m[27]), .Z(pc_a_31__N_1586[25])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i26_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i25_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[26]), .D(branch_target_m[26]), .Z(pc_a_31__N_1586[24])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i25_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i24_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[25]), .D(branch_target_m[25]), .Z(pc_a_31__N_1586[23])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i24_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i23_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[24]), .D(branch_target_m[24]), .Z(pc_a_31__N_1586[22])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i23_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i22_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[23]), .D(branch_target_m[23]), .Z(pc_a_31__N_1586[21])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i22_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i21_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[22]), .D(branch_target_m[22]), .Z(pc_a_31__N_1586[20])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i21_3_lut_4_lut.init = 16'hfb40;
    FD1P3AX wb_data_f_i0_i20 (.D(SHAREDBUS_DAT_O[20]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[20])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i20.GSR = "ENABLED";
    FD1P3AX wb_data_f_i0_i19 (.D(SHAREDBUS_DAT_O[19]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[19])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i19.GSR = "ENABLED";
    LUT4 branch_target_m_31__I_0_i20_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[21]), .D(branch_target_m[21]), .Z(pc_a_31__N_1586[19])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i20_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i19_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[20]), .D(branch_target_m[20]), .Z(pc_a_31__N_1586[18])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i19_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i18_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[19]), .D(branch_target_m[19]), .Z(pc_a_31__N_1586[17])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i18_3_lut_4_lut.init = 16'hfb40;
    FD1P3AX wb_data_f_i0_i18 (.D(SHAREDBUS_DAT_O[18]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[18])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i18.GSR = "ENABLED";
    LUT4 branch_target_m_31__I_0_i17_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[18]), .D(branch_target_m[18]), .Z(pc_a_31__N_1586[16])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i17_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i16_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[17]), .D(branch_target_m[17]), .Z(pc_a_31__N_1586[15])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i16_3_lut_4_lut.init = 16'hfb40;
    FD1P3AX wb_data_f_i0_i17 (.D(SHAREDBUS_DAT_O[17]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[17])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i17.GSR = "ENABLED";
    LUT4 branch_target_m_31__I_0_i15_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[16]), .D(branch_target_m[16]), .Z(pc_a_31__N_1586[14])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i15_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i14_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[15]), .D(branch_target_m[15]), .Z(pc_a_31__N_1586[13])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i14_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i13_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[14]), .D(branch_target_m[14]), .Z(pc_a_31__N_1586[12])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i13_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i12_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[13]), .D(branch_target_m[13]), .Z(pc_a_31__N_1586[11])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i12_3_lut_4_lut.init = 16'hfb40;
    FD1P3AX wb_data_f_i0_i16 (.D(SHAREDBUS_DAT_O[16]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[16])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i16.GSR = "ENABLED";
    LUT4 branch_target_m_31__I_0_i11_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[12]), .D(branch_target_m[12]), .Z(pc_a_31__N_1586[10])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i11_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i10_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[11]), .D(branch_target_m[11]), .Z(pc_a_31__N_1586[9])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i10_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i9_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[10]), .D(branch_target_m[10]), .Z(pc_a_31__N_1586[8])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i9_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i8_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[9]), .D(branch_target_m[9]), .Z(pc_a_31__N_1586[7])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i8_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i7_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[8]), .D(branch_target_m[8]), .Z(pc_a_31__N_1586[6])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i7_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i6_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[7]), .D(branch_target_m[7]), .Z(pc_a_31__N_1586[5])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i6_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i5_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[6]), .D(branch_target_m[6]), .Z(pc_a_31__N_1586[4])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i5_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i4_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[5]), .D(branch_target_m[5]), .Z(pc_a_31__N_1586[3])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i4_3_lut_4_lut.init = 16'hfb40;
    FD1P3AX wb_data_f_i0_i15 (.D(SHAREDBUS_DAT_O[15]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[15])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i15.GSR = "ENABLED";
    LUT4 branch_target_m_31__I_0_i3_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[4]), .D(branch_target_m[4]), .Z(pc_a_31__N_1586[2])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i3_3_lut_4_lut.init = 16'hfb40;
    LUT4 branch_target_m_31__I_0_i2_3_lut_4_lut (.A(n42746), .B(n41459), 
         .C(pc_x[3]), .D(branch_target_m[3]), .Z(pc_a_31__N_1586[1])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_cpu.v(2003[58:81])
    defparam branch_target_m_31__I_0_i2_3_lut_4_lut.init = 16'hfb40;
    FD1P3AX wb_data_f_i0_i14 (.D(SHAREDBUS_DAT_O[14]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[14])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i14.GSR = "ENABLED";
    FD1P3AX wb_data_f_i0_i13 (.D(SHAREDBUS_DAT_O[13]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[13])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i13.GSR = "ENABLED";
    FD1P3AX wb_data_f_i0_i12 (.D(SHAREDBUS_DAT_O[12]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[12])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i12.GSR = "ENABLED";
    LUT4 pc_a_31__I_0_i1_3_lut (.A(pc_a_31__N_1556[0]), .B(pc_a_31__N_1586[0]), 
         .C(branch_taken_m), .Z(pc_a[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i1_3_lut.init = 16'hcaca;
    LUT4 i419_2_lut (.A(i_cyc_o_N_1759), .B(LM32I_CYC_O), .Z(w_clk_cpu_enable_558)) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(829[9] 861[12])
    defparam i419_2_lut.init = 16'h8888;
    FD1P3AX wb_data_f_i0_i11 (.D(SHAREDBUS_DAT_O[11]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[11])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i11.GSR = "ENABLED";
    LUT4 i23410_1_lut (.A(LM32I_CYC_O), .Z(i_cyc_o_N_1754)) /* synthesis lut_function=(!(A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(829[9] 861[12])
    defparam i23410_1_lut.init = 16'h5555;
    FD1P3AX wb_data_f_i0_i10 (.D(SHAREDBUS_DAT_O[10]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[10])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i10.GSR = "ENABLED";
    FD1P3AX wb_data_f_i0_i9 (.D(SHAREDBUS_DAT_O[9]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[9])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i9.GSR = "ENABLED";
    FD1P3AX pc_d_i2_i16 (.D(pc_f[16]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_d[16])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i16.GSR = "ENABLED";
    FD1P3AX wb_data_f_i0_i8 (.D(SHAREDBUS_DAT_O[8]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[8])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i8.GSR = "ENABLED";
    FD1P3AX wb_data_f_i0_i7 (.D(SHAREDBUS_DAT_O[7]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[7])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i7.GSR = "ENABLED";
    CCU2D add_18875_rep_2_15 (.A0(pc_f[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pc_f[16]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n36605), .COUT(n36606), .S0(n22259), .S1(n22258));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_2_15.INIT0 = 16'hfaaa;
    defparam add_18875_rep_2_15.INIT1 = 16'hfaaa;
    defparam add_18875_rep_2_15.INJECT1_0 = "NO";
    defparam add_18875_rep_2_15.INJECT1_1 = "NO";
    FD1P3AX wb_data_f_i0_i6 (.D(SHAREDBUS_DAT_O[6]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[6])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i6.GSR = "ENABLED";
    CCU2D add_18875_rep_2_13 (.A0(pc_f[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pc_f[14]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n36604), .COUT(n36605), .S0(n22261), .S1(n22260));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_2_13.INIT0 = 16'hfaaa;
    defparam add_18875_rep_2_13.INIT1 = 16'hfaaa;
    defparam add_18875_rep_2_13.INJECT1_0 = "NO";
    defparam add_18875_rep_2_13.INJECT1_1 = "NO";
    FD1P3AX wb_data_f_i0_i5 (.D(SHAREDBUS_DAT_O[5]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[5])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i5.GSR = "ENABLED";
    FD1P3AX wb_data_f_i0_i4 (.D(SHAREDBUS_DAT_O[4]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i4.GSR = "ENABLED";
    CCU2D add_18875_rep_2_11 (.A0(pc_f[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pc_f[12]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n36603), .COUT(n36604), .S0(n22263), .S1(n22262));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_2_11.INIT0 = 16'hfaaa;
    defparam add_18875_rep_2_11.INIT1 = 16'hfaaa;
    defparam add_18875_rep_2_11.INJECT1_0 = "NO";
    defparam add_18875_rep_2_11.INJECT1_1 = "NO";
    CCU2D add_18875_rep_2_9 (.A0(pc_f[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pc_f[10]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n36602), .COUT(n36603), .S0(n22265), .S1(n22264));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_2_9.INIT0 = 16'hfaaa;
    defparam add_18875_rep_2_9.INIT1 = 16'hfaaa;
    defparam add_18875_rep_2_9.INJECT1_0 = "NO";
    defparam add_18875_rep_2_9.INJECT1_1 = "NO";
    FD1P3AX wb_data_f_i0_i3 (.D(SHAREDBUS_DAT_O[3]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i3.GSR = "ENABLED";
    FD1P3AX wb_data_f_i0_i2 (.D(SHAREDBUS_DAT_O[2]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i2.GSR = "ENABLED";
    CCU2D add_18875_rep_2_7 (.A0(pc_f[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pc_f[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n36601), .COUT(n36602), .S0(n22267), .S1(n22266));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_2_7.INIT0 = 16'hfaaa;
    defparam add_18875_rep_2_7.INIT1 = 16'hfaaa;
    defparam add_18875_rep_2_7.INJECT1_0 = "NO";
    defparam add_18875_rep_2_7.INJECT1_1 = "NO";
    CCU2D add_18875_rep_2_5 (.A0(pc_f[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pc_f[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n36600), .COUT(n36601), .S0(n22269), .S1(n22268));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_2_5.INIT0 = 16'hfaaa;
    defparam add_18875_rep_2_5.INIT1 = 16'hfaaa;
    defparam add_18875_rep_2_5.INJECT1_0 = "NO";
    defparam add_18875_rep_2_5.INJECT1_1 = "NO";
    FD1P3AX wb_data_f_i0_i1 (.D(SHAREDBUS_DAT_O[1]), .SP(w_clk_cpu_enable_558), 
            .CK(w_clk_cpu), .Q(wb_data_f[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam wb_data_f_i0_i1.GSR = "ENABLED";
    CCU2D add_18875_rep_2_3 (.A0(pc_f[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pc_f[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n36599), .COUT(n36600), .S0(n22271), .S1(n22270));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_2_3.INIT0 = 16'hfaaa;
    defparam add_18875_rep_2_3.INIT1 = 16'hfaaa;
    defparam add_18875_rep_2_3.INJECT1_0 = "NO";
    defparam add_18875_rep_2_3.INJECT1_1 = "NO";
    CCU2D add_18875_rep_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(valid_d), .B1(n41394), .C1(pc_f[2]), .D1(GND_net), 
          .COUT(n36599), .S1(n22272));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_2_1.INIT0 = 16'hF000;
    defparam add_18875_rep_2_1.INIT1 = 16'h8787;
    defparam add_18875_rep_2_1.INJECT1_0 = "NO";
    defparam add_18875_rep_2_1.INJECT1_1 = "NO";
    FD1P3AX i_adr_o__i30 (.D(pc_a[31]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[31] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i30.GSR = "ENABLED";
    FD1P3AX bus_error_f_76 (.D(bus_error_f_N_1764), .SP(w_clk_cpu_enable_587), 
            .CK(w_clk_cpu), .Q(bus_error_f)) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam bus_error_f_76.GSR = "ENABLED";
    FD1P3AX i_adr_o__i29 (.D(pc_a[30]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[30] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i29.GSR = "ENABLED";
    CCU2D add_18875_rep_3_31 (.A0(n22244), .B0(n41375), .C0(\branch_target_d[30] ), 
          .D0(GND_net), .A1(n22243), .B1(n41375), .C1(\branch_target_d[31] ), 
          .D1(GND_net), .CIN(n36597), .S0(pc_a_31__N_1556[28]), .S1(pc_a_31__N_1556[29]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_3_31.INIT0 = 16'hd2e2;
    defparam add_18875_rep_3_31.INIT1 = 16'hd2e2;
    defparam add_18875_rep_3_31.INJECT1_0 = "NO";
    defparam add_18875_rep_3_31.INJECT1_1 = "NO";
    FD1P3AX i_adr_o__i28 (.D(pc_a[29]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[29] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i28.GSR = "ENABLED";
    CCU2D add_18875_rep_3_29 (.A0(n22246), .B0(n41375), .C0(\branch_target_d[28] ), 
          .D0(GND_net), .A1(n22245), .B1(n41375), .C1(\branch_target_d[29] ), 
          .D1(GND_net), .CIN(n36596), .COUT(n36597), .S0(pc_a_31__N_1556[26]), 
          .S1(pc_a_31__N_1556[27]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_3_29.INIT0 = 16'hd2e2;
    defparam add_18875_rep_3_29.INIT1 = 16'hd2e2;
    defparam add_18875_rep_3_29.INJECT1_0 = "NO";
    defparam add_18875_rep_3_29.INJECT1_1 = "NO";
    FD1P3AX i_adr_o__i27 (.D(pc_a[28]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[28] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i27.GSR = "ENABLED";
    CCU2D add_18875_rep_3_27 (.A0(n22248), .B0(n41375), .C0(\branch_target_d[26] ), 
          .D0(GND_net), .A1(n22247), .B1(n41375), .C1(\branch_target_d[27] ), 
          .D1(GND_net), .CIN(n36595), .COUT(n36596), .S0(pc_a_31__N_1556[24]), 
          .S1(pc_a_31__N_1556[25]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_3_27.INIT0 = 16'hd2e2;
    defparam add_18875_rep_3_27.INIT1 = 16'hd2e2;
    defparam add_18875_rep_3_27.INJECT1_0 = "NO";
    defparam add_18875_rep_3_27.INJECT1_1 = "NO";
    FD1P3AX i_adr_o__i26 (.D(pc_a[27]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[27] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i26.GSR = "ENABLED";
    CCU2D add_18875_rep_3_25 (.A0(n22250), .B0(n41375), .C0(\branch_target_d[24] ), 
          .D0(GND_net), .A1(n22249), .B1(n41375), .C1(\branch_target_d[25] ), 
          .D1(GND_net), .CIN(n36594), .COUT(n36595), .S0(pc_a_31__N_1556[22]), 
          .S1(pc_a_31__N_1556[23]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_3_25.INIT0 = 16'hd2e2;
    defparam add_18875_rep_3_25.INIT1 = 16'hd2e2;
    defparam add_18875_rep_3_25.INJECT1_0 = "NO";
    defparam add_18875_rep_3_25.INJECT1_1 = "NO";
    FD1P3AX i_adr_o__i25 (.D(pc_a[26]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[26] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i25.GSR = "ENABLED";
    FD1P3AX i_adr_o__i24 (.D(pc_a[25]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[25] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i24.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i31 (.D(pc_a[31]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_f[31])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i31.GSR = "ENABLED";
    CCU2D add_18875_rep_3_23 (.A0(n22252), .B0(n41375), .C0(\branch_target_d[22] ), 
          .D0(GND_net), .A1(n22251), .B1(n41375), .C1(\branch_target_d[23] ), 
          .D1(GND_net), .CIN(n36593), .COUT(n36594), .S0(pc_a_31__N_1556[20]), 
          .S1(pc_a_31__N_1556[21]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_3_23.INIT0 = 16'hd2e2;
    defparam add_18875_rep_3_23.INIT1 = 16'hd2e2;
    defparam add_18875_rep_3_23.INJECT1_0 = "NO";
    defparam add_18875_rep_3_23.INJECT1_1 = "NO";
    CCU2D add_18875_rep_3_21 (.A0(n22254), .B0(n41375), .C0(\branch_target_d[20] ), 
          .D0(GND_net), .A1(n22253), .B1(n41375), .C1(\branch_target_d[21] ), 
          .D1(GND_net), .CIN(n36592), .COUT(n36593), .S0(pc_a_31__N_1556[18]), 
          .S1(pc_a_31__N_1556[19]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_3_21.INIT0 = 16'hd2e2;
    defparam add_18875_rep_3_21.INIT1 = 16'hd2e2;
    defparam add_18875_rep_3_21.INJECT1_0 = "NO";
    defparam add_18875_rep_3_21.INJECT1_1 = "NO";
    FD1P3AX i_adr_o__i23 (.D(pc_a[24]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[24] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i23.GSR = "ENABLED";
    FD1P3AX i_adr_o__i22 (.D(pc_a[23]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[23] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i22.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i30 (.D(pc_a[30]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_f[30])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i30.GSR = "ENABLED";
    CCU2D add_18875_rep_3_19 (.A0(n22256), .B0(n41375), .C0(\branch_target_d[18] ), 
          .D0(GND_net), .A1(n22255), .B1(n41375), .C1(\branch_target_d[19] ), 
          .D1(GND_net), .CIN(n36591), .COUT(n36592), .S0(pc_a_31__N_1556[16]), 
          .S1(pc_a_31__N_1556[17]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_3_19.INIT0 = 16'hd2e2;
    defparam add_18875_rep_3_19.INIT1 = 16'hd2e2;
    defparam add_18875_rep_3_19.INJECT1_0 = "NO";
    defparam add_18875_rep_3_19.INJECT1_1 = "NO";
    CCU2D add_18875_rep_3_17 (.A0(n22258), .B0(n41375), .C0(\branch_target_d[16] ), 
          .D0(GND_net), .A1(n22257), .B1(n41375), .C1(\branch_target_d[17] ), 
          .D1(GND_net), .CIN(n36590), .COUT(n36591), .S0(pc_a_31__N_1556[14]), 
          .S1(pc_a_31__N_1556[15]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_3_17.INIT0 = 16'hd2e2;
    defparam add_18875_rep_3_17.INIT1 = 16'hd2e2;
    defparam add_18875_rep_3_17.INJECT1_0 = "NO";
    defparam add_18875_rep_3_17.INJECT1_1 = "NO";
    FD1P3AX i_adr_o__i21 (.D(pc_a[22]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[22] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i21.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i29 (.D(pc_a[29]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_f[29])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i29.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i28 (.D(pc_a[28]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_f[28])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i28.GSR = "ENABLED";
    CCU2D add_18875_rep_3_15 (.A0(n22260), .B0(n41375), .C0(\branch_target_d[14] ), 
          .D0(GND_net), .A1(n22259), .B1(n41375), .C1(\branch_target_d[15] ), 
          .D1(GND_net), .CIN(n36589), .COUT(n36590), .S0(pc_a_31__N_1556[12]), 
          .S1(pc_a_31__N_1556[13]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_3_15.INIT0 = 16'hd2e2;
    defparam add_18875_rep_3_15.INIT1 = 16'hd2e2;
    defparam add_18875_rep_3_15.INJECT1_0 = "NO";
    defparam add_18875_rep_3_15.INJECT1_1 = "NO";
    FD1P3AX i_adr_o__i20 (.D(pc_a[21]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[21] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i20.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i27 (.D(pc_a[27]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_f[27])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i27.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i26 (.D(pc_a[26]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_f[26])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i26.GSR = "ENABLED";
    CCU2D add_18875_rep_3_13 (.A0(n22262), .B0(n41375), .C0(\branch_target_d[12] ), 
          .D0(GND_net), .A1(n22261), .B1(n41375), .C1(\branch_target_d[13] ), 
          .D1(GND_net), .CIN(n36588), .COUT(n36589), .S0(pc_a_31__N_1556[10]), 
          .S1(pc_a_31__N_1556[11]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_3_13.INIT0 = 16'hd2e2;
    defparam add_18875_rep_3_13.INIT1 = 16'hd2e2;
    defparam add_18875_rep_3_13.INJECT1_0 = "NO";
    defparam add_18875_rep_3_13.INJECT1_1 = "NO";
    FD1P3AX i_adr_o__i19 (.D(pc_a[20]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[20] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i19.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i25 (.D(pc_a[25]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_f[25])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i25.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i24 (.D(pc_a[24]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_f[24])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i24.GSR = "ENABLED";
    FD1P3AX i_adr_o__i18 (.D(pc_a[19]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[19] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i18.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i23 (.D(pc_a[23]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_f[23])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i23.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i22 (.D(pc_a[22]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_f[22])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i22.GSR = "ENABLED";
    FD1P3AX i_adr_o__i17 (.D(pc_a[18]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[18] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i17.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i21 (.D(pc_a[21]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_f[21])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i21.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i20 (.D(pc_a[20]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_f[20])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i20.GSR = "ENABLED";
    FD1P3AX i_adr_o__i16 (.D(pc_a[17]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[17] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i16.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i19 (.D(pc_a[19]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_f[19])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i19.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i18 (.D(pc_a[18]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_f[18])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i18.GSR = "ENABLED";
    CCU2D add_18875_rep_3_7 (.A0(n22268), .B0(n41375), .C0(\branch_target_d[6] ), 
          .D0(GND_net), .A1(n22267), .B1(n41375), .C1(\branch_target_d[7] ), 
          .D1(GND_net), .CIN(n36585), .COUT(n36586), .S0(pc_a_31__N_1556[4]), 
          .S1(pc_a_31__N_1556[5]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_3_7.INIT0 = 16'hd2e2;
    defparam add_18875_rep_3_7.INIT1 = 16'hd2e2;
    defparam add_18875_rep_3_7.INJECT1_0 = "NO";
    defparam add_18875_rep_3_7.INJECT1_1 = "NO";
    FD1P3AX i_adr_o__i15 (.D(pc_a[16]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[16] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i15.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i17 (.D(pc_a[17]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_f[17])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i17.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i16 (.D(pc_a[16]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_f[16])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i16.GSR = "ENABLED";
    CCU2D add_18875_rep_2_31 (.A0(pc_f[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n36613), .S0(n22243));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_2_31.INIT0 = 16'hfaaa;
    defparam add_18875_rep_2_31.INIT1 = 16'h0000;
    defparam add_18875_rep_2_31.INJECT1_0 = "NO";
    defparam add_18875_rep_2_31.INJECT1_1 = "NO";
    CCU2D add_18875_rep_2_29 (.A0(pc_f[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pc_f[30]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n36612), .COUT(n36613), .S0(n22245), .S1(n22244));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_2_29.INIT0 = 16'hfaaa;
    defparam add_18875_rep_2_29.INIT1 = 16'hfaaa;
    defparam add_18875_rep_2_29.INJECT1_0 = "NO";
    defparam add_18875_rep_2_29.INJECT1_1 = "NO";
    CCU2D add_18875_rep_2_27 (.A0(pc_f[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pc_f[28]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n36611), .COUT(n36612), .S0(n22247), .S1(n22246));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_2_27.INIT0 = 16'hfaaa;
    defparam add_18875_rep_2_27.INIT1 = 16'hfaaa;
    defparam add_18875_rep_2_27.INJECT1_0 = "NO";
    defparam add_18875_rep_2_27.INJECT1_1 = "NO";
    CCU2D add_18875_rep_2_25 (.A0(pc_f[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pc_f[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n36610), .COUT(n36611), .S0(n22249), .S1(n22248));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_2_25.INIT0 = 16'hfaaa;
    defparam add_18875_rep_2_25.INIT1 = 16'hfaaa;
    defparam add_18875_rep_2_25.INJECT1_0 = "NO";
    defparam add_18875_rep_2_25.INJECT1_1 = "NO";
    CCU2D add_18875_rep_2_23 (.A0(pc_f[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pc_f[24]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n36609), .COUT(n36610), .S0(n22251), .S1(n22250));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_2_23.INIT0 = 16'hfaaa;
    defparam add_18875_rep_2_23.INIT1 = 16'hfaaa;
    defparam add_18875_rep_2_23.INJECT1_0 = "NO";
    defparam add_18875_rep_2_23.INJECT1_1 = "NO";
    FD1P3AX pc_d_i2_i15 (.D(pc_f[15]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_d[15])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_d_i2_i15.GSR = "ENABLED";
    FD1P3AX i_adr_o__i14 (.D(pc_a[15]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[15] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i14.GSR = "ENABLED";
    FD1P3AX i_adr_o__i13 (.D(pc_a[14]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[14] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i13.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i15 (.D(pc_a[15]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_f[15])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i15.GSR = "ENABLED";
    CCU2D add_18875_rep_3_9 (.A0(n22266), .B0(n41375), .C0(\branch_target_d[8] ), 
          .D0(GND_net), .A1(n22265), .B1(n41375), .C1(\branch_target_d[9] ), 
          .D1(GND_net), .CIN(n36586), .COUT(n36587), .S0(pc_a_31__N_1556[6]), 
          .S1(pc_a_31__N_1556[7]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_3_9.INIT0 = 16'hd2e2;
    defparam add_18875_rep_3_9.INIT1 = 16'hd2e2;
    defparam add_18875_rep_3_9.INJECT1_0 = "NO";
    defparam add_18875_rep_3_9.INJECT1_1 = "NO";
    FD1P3AX i_adr_o__i12 (.D(pc_a[13]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[13] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i12.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i14 (.D(pc_a[14]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_f[14])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i14.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i13 (.D(pc_a[13]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_f[13])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i13.GSR = "ENABLED";
    CCU2D add_18875_rep_3_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(valid_d), .B1(n41394), .C1(GND_net), .D1(GND_net), 
          .COUT(n36583));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_3_1.INIT0 = 16'hF000;
    defparam add_18875_rep_3_1.INIT1 = 16'hffff;
    defparam add_18875_rep_3_1.INJECT1_0 = "NO";
    defparam add_18875_rep_3_1.INJECT1_1 = "NO";
    CCU2D add_18875_rep_2_21 (.A0(pc_f[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(pc_f[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n36608), .COUT(n36609), .S0(n22253), .S1(n22252));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_2_21.INIT0 = 16'hfaaa;
    defparam add_18875_rep_2_21.INIT1 = 16'hfaaa;
    defparam add_18875_rep_2_21.INJECT1_0 = "NO";
    defparam add_18875_rep_2_21.INJECT1_1 = "NO";
    FD1P3AX i_adr_o__i11 (.D(pc_a[12]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[12] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i11.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i12 (.D(pc_a[12]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_f[12])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i12.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i11 (.D(pc_a[11]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_f[11])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i11.GSR = "ENABLED";
    CCU2D add_18875_rep_3_5 (.A0(n22270), .B0(n41375), .C0(\branch_target_d[4] ), 
          .D0(GND_net), .A1(n22269), .B1(n41375), .C1(\branch_target_d[5] ), 
          .D1(GND_net), .CIN(n36584), .COUT(n36585), .S0(pc_a_31__N_1556[2]), 
          .S1(pc_a_31__N_1556[3]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_3_5.INIT0 = 16'hd2e2;
    defparam add_18875_rep_3_5.INIT1 = 16'hd2e2;
    defparam add_18875_rep_3_5.INJECT1_0 = "NO";
    defparam add_18875_rep_3_5.INJECT1_1 = "NO";
    FD1P3AX i_adr_o__i10 (.D(pc_a[11]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[11] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i10.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i10 (.D(pc_a[10]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_f[10])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i10.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i9 (.D(pc_a[9]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_f[9])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i9.GSR = "ENABLED";
    CCU2D add_18875_rep_3_11 (.A0(n22264), .B0(n41375), .C0(\branch_target_d[10] ), 
          .D0(GND_net), .A1(n22263), .B1(n41375), .C1(\branch_target_d[11] ), 
          .D1(GND_net), .CIN(n36587), .COUT(n36588), .S0(pc_a_31__N_1556[8]), 
          .S1(pc_a_31__N_1556[9]));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(511[6:25])
    defparam add_18875_rep_3_11.INIT0 = 16'hd2e2;
    defparam add_18875_rep_3_11.INIT1 = 16'hd2e2;
    defparam add_18875_rep_3_11.INJECT1_0 = "NO";
    defparam add_18875_rep_3_11.INJECT1_1 = "NO";
    FD1P3AX i_adr_o__i9 (.D(pc_a[10]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[10] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i9.GSR = "ENABLED";
    FD1P3AX i_adr_o__i8 (.D(pc_a[9]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[9] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i8.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i8 (.D(pc_a[8]), .SP(w_clk_cpu_enable_983), .CK(w_clk_cpu), 
            .Q(pc_f[8])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i8.GSR = "ENABLED";
    FD1P3AX i_adr_o__i7 (.D(pc_a[8]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[8] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i7.GSR = "ENABLED";
    FD1P3AX i_adr_o__i6 (.D(pc_a[7]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[7] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i6.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i7 (.D(pc_a[7]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_f[7])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i7.GSR = "ENABLED";
    FD1P3AX i_adr_o__i5 (.D(pc_a[6]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[6] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i5.GSR = "ENABLED";
    FD1P3AX i_adr_o__i4 (.D(pc_a[5]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[5] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i4.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i6 (.D(pc_a[6]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_f[6])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i6.GSR = "ENABLED";
    FD1P3AX i_adr_o__i3 (.D(pc_a[4]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[4] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i3.GSR = "ENABLED";
    FD1P3AX i_adr_o__i2 (.D(pc_a[3]), .SP(w_clk_cpu_enable_763), .CK(w_clk_cpu), 
            .Q(\LM32I_ADR_O[3] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(807[5] 862[8])
    defparam i_adr_o__i2.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i5 (.D(pc_a[5]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_f[5])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i5.GSR = "ENABLED";
    LUT4 i12_4_lut (.A(n42740), .B(n41479), .C(LM32I_CYC_O), .D(n38871), 
         .Z(w_clk_cpu_enable_587)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam i12_4_lut.init = 16'hca0a;
    FD1P3AX pc_m_i2_i31 (.D(pc_x[31]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[31])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i31.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i30 (.D(pc_x[30]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[30])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i30.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i4 (.D(pc_a[4]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_f[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i4.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i29 (.D(pc_x[29]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[29])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i29.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i28 (.D(pc_x[28]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[28])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i28.GSR = "ENABLED";
    FD1P3AY pc_f_i2_i3 (.D(pc_a[3]), .SP(w_clk_cpu_enable_914), .CK(w_clk_cpu), 
            .Q(pc_f[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_f_i2_i3.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i27 (.D(pc_x[27]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[27])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i27.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i26 (.D(pc_x[26]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[26])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i26.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i25 (.D(pc_x[25]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[25])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i25.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i24 (.D(pc_x[24]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[24])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i24.GSR = "ENABLED";
    FD1P3AX bus_error_d_78 (.D(bus_error_f), .SP(w_clk_cpu_enable_914), 
            .CK(w_clk_cpu), .Q(bus_error_d));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam bus_error_d_78.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i23 (.D(pc_x[23]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[23])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i23.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i22 (.D(pc_x[22]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[22])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i22.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i31 (.D(wb_data_f[31]), .SP(w_clk_cpu_enable_914), 
            .CK(w_clk_cpu), .Q(\instruction_d[31] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i31.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i21 (.D(pc_x[21]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[21])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i21.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i20 (.D(pc_x[20]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[20])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i20.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i30 (.D(wb_data_f[30]), .SP(w_clk_cpu_enable_914), 
            .CK(w_clk_cpu), .Q(\instruction_d[30] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i30.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i19 (.D(pc_x[19]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[19])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i19.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i18 (.D(pc_x[18]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[18])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i18.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i29 (.D(wb_data_f[29]), .SP(w_clk_cpu_enable_914), 
            .CK(w_clk_cpu), .Q(\logic_op_d[3] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i29.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i17 (.D(pc_x[17]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[17])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i17.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i16 (.D(pc_x[16]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[16])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i16.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i28 (.D(wb_data_f[28]), .SP(w_clk_cpu_enable_914), 
            .CK(w_clk_cpu), .Q(sign_extend_d)) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i28.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i15 (.D(pc_x[15]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[15])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i15.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i14 (.D(pc_x[14]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[14])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i14.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i27 (.D(wb_data_f[27]), .SP(w_clk_cpu_enable_914), 
            .CK(w_clk_cpu), .Q(size_d[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i27.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i13 (.D(pc_x[13]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[13])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i13.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i12 (.D(pc_x[12]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[12])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i12.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i26 (.D(wb_data_f[26]), .SP(w_clk_cpu_enable_983), 
            .CK(w_clk_cpu), .Q(size_d[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i26.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i11 (.D(pc_x[11]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[11])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i11.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i10 (.D(pc_x[10]), .SP(w_clk_cpu_enable_878), .CK(w_clk_cpu), 
            .Q(pc_m[10])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i10.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i25 (.D(wb_data_f[25]), .SP(w_clk_cpu_enable_914), 
            .CK(w_clk_cpu), .Q(read_idx_0_d[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i25.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i9 (.D(pc_x[9]), .SP(w_clk_cpu_enable_985), .CK(w_clk_cpu), 
            .Q(pc_m[9])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i9.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i8 (.D(pc_x[8]), .SP(w_clk_cpu_enable_985), .CK(w_clk_cpu), 
            .Q(pc_m[8])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i8.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i24 (.D(wb_data_f[24]), .SP(w_clk_cpu_enable_914), 
            .CK(w_clk_cpu), .Q(read_idx_0_d[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i24.GSR = "ENABLED";
    LUT4 pc_a_31__I_0_i30_3_lut (.A(pc_a_31__N_1556[29]), .B(pc_a_31__N_1586[29]), 
         .C(branch_taken_m), .Z(pc_a[31])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(503[2] 511[25])
    defparam pc_a_31__I_0_i30_3_lut.init = 16'hcaca;
    FD1P3AX pc_m_i2_i7 (.D(pc_x[7]), .SP(w_clk_cpu_enable_985), .CK(w_clk_cpu), 
            .Q(pc_m[7])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i7.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i6 (.D(pc_x[6]), .SP(w_clk_cpu_enable_985), .CK(w_clk_cpu), 
            .Q(pc_m[6])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i6.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i23 (.D(wb_data_f[23]), .SP(w_clk_cpu_enable_914), 
            .CK(w_clk_cpu), .Q(read_idx_0_d[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i23.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i5 (.D(pc_x[5]), .SP(w_clk_cpu_enable_985), .CK(w_clk_cpu), 
            .Q(pc_m[5])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i5.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i4 (.D(pc_x[4]), .SP(w_clk_cpu_enable_985), .CK(w_clk_cpu), 
            .Q(pc_m[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i4.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i22 (.D(wb_data_f[22]), .SP(w_clk_cpu_enable_914), 
            .CK(w_clk_cpu), .Q(read_idx_0_d[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i22.GSR = "ENABLED";
    FD1P3AX pc_m_i2_i3 (.D(pc_x[3]), .SP(w_clk_cpu_enable_985), .CK(w_clk_cpu), 
            .Q(pc_m[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_m_i2_i3.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i31 (.D(pc_d[31]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[31])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i31.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i21 (.D(wb_data_f[21]), .SP(w_clk_cpu_enable_914), 
            .CK(w_clk_cpu), .Q(read_idx_0_d[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i21.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i30 (.D(pc_d[30]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[30])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i30.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i29 (.D(pc_d[29]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[29])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i29.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i20 (.D(wb_data_f[20]), .SP(w_clk_cpu_enable_983), 
            .CK(w_clk_cpu), .Q(read_idx_1_d[4])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i20.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i28 (.D(pc_d[28]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[28])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i28.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i27 (.D(pc_d[27]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[27])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i27.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i19 (.D(wb_data_f[19]), .SP(w_clk_cpu_enable_983), 
            .CK(w_clk_cpu), .Q(read_idx_1_d[3])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i19.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i26 (.D(pc_d[26]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[26])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i26.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i25 (.D(pc_d[25]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[25])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i25.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i18 (.D(wb_data_f[18]), .SP(w_clk_cpu_enable_983), 
            .CK(w_clk_cpu), .Q(read_idx_1_d[2])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i18.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i24 (.D(pc_d[24]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[24])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i24.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i23 (.D(pc_d[23]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[23])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i23.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i17 (.D(wb_data_f[17]), .SP(w_clk_cpu_enable_983), 
            .CK(w_clk_cpu), .Q(read_idx_1_d[1])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i17.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i22 (.D(pc_d[22]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[22])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i22.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i21 (.D(pc_d[21]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[21])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i21.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i16 (.D(wb_data_f[16]), .SP(w_clk_cpu_enable_983), 
            .CK(w_clk_cpu), .Q(read_idx_1_d[0])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i16.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i20 (.D(pc_d[20]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[20])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i20.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i19 (.D(pc_d[19]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[19])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i19.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i15 (.D(wb_data_f[15]), .SP(w_clk_cpu_enable_983), 
            .CK(w_clk_cpu), .Q(\instruction_d[15] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i15.GSR = "ENABLED";
    FD1P3AX pc_x_i2_i18 (.D(pc_d[18]), .SP(w_clk_cpu_enable_984), .CK(w_clk_cpu), 
            .Q(pc_x[18])) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(605[8] 615[11])
    defparam pc_x_i2_i18.GSR = "ENABLED";
    FD1P3AX instruction_d_i0_i14 (.D(wb_data_f[14]), .SP(w_clk_cpu_enable_983), 
            .CK(w_clk_cpu), .Q(\instruction_d[14] )) /* synthesis LSE_LINE_FILE_ID=21, LSE_LCOL=5, LSE_RCOL=6, LSE_LLINE=804, LSE_RLINE=896 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_instruction_unit.v(878[5] 886[8])
    defparam instruction_d_i0_i14.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \lm32_debug(watchpoints=32'b0) 
//

module \lm32_debug(watchpoints=32'b0)  (dc_re, w_clk_cpu, dc_re_N_2934, 
            \operand_1_x[1] ) /* synthesis syn_module_defined=1 */ ;
    output dc_re;
    input w_clk_cpu;
    input dc_re_N_2934;
    input \operand_1_x[1] ;
    
    wire w_clk_cpu /* synthesis SET_AS_NETWORK=w_clk_cpu, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(22[6:15])
    
    FD1P3AX dc_re_10 (.D(\operand_1_x[1] ), .SP(dc_re_N_2934), .CK(w_clk_cpu), 
            .Q(dc_re));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_debug.v(296[5] 299[8])
    defparam dc_re_10.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module lm32_decoder
//

module lm32_decoder (size_d, sign_extend_d, \instruction_d[30] , \instruction_d[31] , 
            \logic_op_d[3] , x_result_sel_csr_d, \instruction_d[0] , n1792, 
            \instruction_d[15] , n1777, n41397, \instruction_d[7] , 
            n1785, \instruction_d[6] , n1786, \instruction_d[5] , n1787, 
            \instruction_d[4] , n1788, \instruction_d[3] , n1789, \instruction_d[2] , 
            n1790, \instruction_d[1] , n1791, n41419, n41376, adder_op_d_N_1339, 
            n41361, n41364, n42740, cycles_5__N_2495, n41345, n13, 
            w_clk_cpu_enable_958, n18875, x_result_sel_sext_N_1782, x_bypass_enable_d, 
            m_bypass_enable_d, read_idx_0_d, eret_d, bret_d, sign_extend_immediate, 
            bus_error_d, n41199, n41367, n41417, n22236, \instruction_d[12] , 
            n2, n2_adj_3, n2_adj_4, n2_adj_5, n2_adj_6, n2_adj_7, 
            n2_adj_8, n2_adj_9, \instruction_d[8] , n2_adj_10, \instruction_d[9] , 
            n2_adj_11, \instruction_d[10] , n2_adj_12, pc_f, \bypass_data_0[31] , 
            \d_result_0[31] , \bypass_data_0[30] , \d_result_0[30] , \bypass_data_0[29] , 
            \d_result_0[29] , \bypass_data_0[28] , \d_result_0[28] , \bypass_data_0[27] , 
            \d_result_0[27] , n2_adj_13, \bypass_data_0[26] , \d_result_0[26] , 
            \bypass_data_0[25] , \d_result_0[25] , \bypass_data_0[24] , 
            \d_result_0[24] , \bypass_data_0[23] , \d_result_0[23] , n22224, 
            \instruction_d[11] , n2_adj_14, \bypass_data_0[22] , \d_result_0[22] , 
            \bypass_data_0[21] , \d_result_0[21] , \bypass_data_0[20] , 
            \d_result_0[20] , \bypass_data_0[19] , \d_result_0[19] , \bypass_data_0[18] , 
            \d_result_0[18] , \bypass_data_0[17] , \d_result_0[17] , \bypass_data_0[16] , 
            \d_result_0[16] , \bypass_data_0[15] , \d_result_0[15] , \bypass_data_0[14] , 
            \d_result_0[14] , \bypass_data_0[13] , \d_result_0[13] , \bypass_data_0[12] , 
            \d_result_0[12] , \bypass_data_0[11] , \d_result_0[11] , \bypass_data_0[10] , 
            \d_result_0[10] , \bypass_data_0[9] , \d_result_0[9] , n42722, 
            \bypass_data_0[8] , \d_result_0[8] , \bypass_data_0[7] , \d_result_0[7] , 
            \bypass_data_0[6] , \d_result_0[6] , n41384, \bypass_data_0[5] , 
            \d_result_0[5] , \bypass_data_0[4] , \d_result_0[4] , n2_adj_15, 
            \bypass_data_0[3] , \d_result_0[3] , \instruction_d[14] , 
            n2_adj_16, \bypass_data_0[2] , \d_result_0[2] , \instruction_d[13] , 
            n2_adj_17, n41407, n1765, n1762, n1763, n1766, n1767, 
            n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, 
            n1776, n1764, read_idx_1_d, \write_idx_4__N_1770[1] , bypass_data_1, 
            n1, n1_adj_18, n1_adj_19, n41394, n1_adj_20, n1_adj_21, 
            n1_adj_22, n1_adj_23, n1_adj_24, n1_adj_25, n1_adj_26, 
            n1_adj_27, n1_adj_28, n1_adj_29, n1_adj_30, n1_adj_31, 
            n1_adj_32, n1_adj_33, branch_d, n1_adj_34, n1_adj_35, 
            n1_adj_36, n1_adj_37, n1_adj_38, n1_adj_39, n1_adj_40, 
            n1_adj_41, n1_adj_42, n1_adj_43, n1_adj_44, n41466, x_result_sel_add_N_1785, 
            n1_adj_45, n1_adj_46, n1_adj_47, n1_adj_48, raw_x_1, raw_x_0, 
            interlock_N_1327, n41411, raw_m_0, interlock_N_1333, n41406, 
            store_d, write_enable_N_1809, w_result_sel_mul_d, n25722, 
            scall_d, break_d, \write_idx_d[4] , \write_idx_d[3] , \write_idx_d[2] , 
            n25724, n41380, \write_idx_d[0] , branch_predict_d, m_result_sel_shift_d) /* synthesis syn_module_defined=1 */ ;
    input [1:0]size_d;
    input sign_extend_d;
    input \instruction_d[30] ;
    input \instruction_d[31] ;
    input \logic_op_d[3] ;
    output x_result_sel_csr_d;
    input \instruction_d[0] ;
    output n1792;
    input \instruction_d[15] ;
    output n1777;
    output n41397;
    input \instruction_d[7] ;
    output n1785;
    input \instruction_d[6] ;
    output n1786;
    input \instruction_d[5] ;
    output n1787;
    input \instruction_d[4] ;
    output n1788;
    input \instruction_d[3] ;
    output n1789;
    input \instruction_d[2] ;
    output n1790;
    input \instruction_d[1] ;
    output n1791;
    output n41419;
    output n41376;
    output adder_op_d_N_1339;
    output n41361;
    output n41364;
    input n42740;
    input cycles_5__N_2495;
    output n41345;
    input n13;
    input w_clk_cpu_enable_958;
    output n18875;
    output x_result_sel_sext_N_1782;
    output x_bypass_enable_d;
    output m_bypass_enable_d;
    input [4:0]read_idx_0_d;
    output eret_d;
    output bret_d;
    output sign_extend_immediate;
    input bus_error_d;
    output n41199;
    output n41367;
    output n41417;
    output n22236;
    input \instruction_d[12] ;
    output n2;
    output n2_adj_3;
    output n2_adj_4;
    output n2_adj_5;
    output n2_adj_6;
    output n2_adj_7;
    output n2_adj_8;
    output n2_adj_9;
    input \instruction_d[8] ;
    output n2_adj_10;
    input \instruction_d[9] ;
    output n2_adj_11;
    input \instruction_d[10] ;
    output n2_adj_12;
    input [31:2]pc_f;
    input \bypass_data_0[31] ;
    output \d_result_0[31] ;
    input \bypass_data_0[30] ;
    output \d_result_0[30] ;
    input \bypass_data_0[29] ;
    output \d_result_0[29] ;
    input \bypass_data_0[28] ;
    output \d_result_0[28] ;
    input \bypass_data_0[27] ;
    output \d_result_0[27] ;
    output n2_adj_13;
    input \bypass_data_0[26] ;
    output \d_result_0[26] ;
    input \bypass_data_0[25] ;
    output \d_result_0[25] ;
    input \bypass_data_0[24] ;
    output \d_result_0[24] ;
    input \bypass_data_0[23] ;
    output \d_result_0[23] ;
    output n22224;
    input \instruction_d[11] ;
    output n2_adj_14;
    input \bypass_data_0[22] ;
    output \d_result_0[22] ;
    input \bypass_data_0[21] ;
    output \d_result_0[21] ;
    input \bypass_data_0[20] ;
    output \d_result_0[20] ;
    input \bypass_data_0[19] ;
    output \d_result_0[19] ;
    input \bypass_data_0[18] ;
    output \d_result_0[18] ;
    input \bypass_data_0[17] ;
    output \d_result_0[17] ;
    input \bypass_data_0[16] ;
    output \d_result_0[16] ;
    input \bypass_data_0[15] ;
    output \d_result_0[15] ;
    input \bypass_data_0[14] ;
    output \d_result_0[14] ;
    input \bypass_data_0[13] ;
    output \d_result_0[13] ;
    input \bypass_data_0[12] ;
    output \d_result_0[12] ;
    input \bypass_data_0[11] ;
    output \d_result_0[11] ;
    input \bypass_data_0[10] ;
    output \d_result_0[10] ;
    input \bypass_data_0[9] ;
    output \d_result_0[9] ;
    output n42722;
    input \bypass_data_0[8] ;
    output \d_result_0[8] ;
    input \bypass_data_0[7] ;
    output \d_result_0[7] ;
    input \bypass_data_0[6] ;
    output \d_result_0[6] ;
    output n41384;
    input \bypass_data_0[5] ;
    output \d_result_0[5] ;
    input \bypass_data_0[4] ;
    output \d_result_0[4] ;
    output n2_adj_15;
    input \bypass_data_0[3] ;
    output \d_result_0[3] ;
    input \instruction_d[14] ;
    output n2_adj_16;
    input \bypass_data_0[2] ;
    output \d_result_0[2] ;
    input \instruction_d[13] ;
    output n2_adj_17;
    output n41407;
    output n1765;
    output n1762;
    output n1763;
    output n1766;
    output n1767;
    output n1768;
    output n1769;
    output n1770;
    output n1771;
    output n1772;
    output n1773;
    output n1774;
    output n1775;
    output n1776;
    output n1764;
    input [4:0]read_idx_1_d;
    output \write_idx_4__N_1770[1] ;
    input [31:0]bypass_data_1;
    output n1;
    output n1_adj_18;
    output n1_adj_19;
    output n41394;
    output n1_adj_20;
    output n1_adj_21;
    output n1_adj_22;
    output n1_adj_23;
    output n1_adj_24;
    output n1_adj_25;
    output n1_adj_26;
    output n1_adj_27;
    output n1_adj_28;
    output n1_adj_29;
    output n1_adj_30;
    output n1_adj_31;
    output n1_adj_32;
    output n1_adj_33;
    output branch_d;
    output n1_adj_34;
    output n1_adj_35;
    output n1_adj_36;
    output n1_adj_37;
    output n1_adj_38;
    output n1_adj_39;
    output n1_adj_40;
    output n1_adj_41;
    output n1_adj_42;
    output n1_adj_43;
    output n1_adj_44;
    output n41466;
    output x_result_sel_add_N_1785;
    output n1_adj_45;
    output n1_adj_46;
    output n1_adj_47;
    output n1_adj_48;
    input raw_x_1;
    input raw_x_0;
    output interlock_N_1327;
    input n41411;
    input raw_m_0;
    output interlock_N_1333;
    output n41406;
    output store_d;
    output write_enable_N_1809;
    output w_result_sel_mul_d;
    output n25722;
    output scall_d;
    output break_d;
    output \write_idx_d[4] ;
    output \write_idx_d[3] ;
    output \write_idx_d[2] ;
    output n25724;
    output n41380;
    output \write_idx_d[0] ;
    output branch_predict_d;
    output m_result_sel_shift_d;
    
    
    wire n23666, n41515, n41463, n41499, n41427, n41533, n41437, 
        n41436, n41434, bra, n41527, n39110, n41528, n41464, n41439, 
        n39002, n41538, n41460, n41396, n41532, n41446, n41433, 
        n8, n38976, n7, n40446, n32034, n39220, n31609, n39191, 
        n58, n8_adj_3651, n23, n41312, n39162, n41494, n10, n40445, 
        n40444, n39005, n20, n6, n41558, n41559, n41486, n41485, 
        n41477, n41631, n39042, n40091, n41138, n41137, n41139, 
        n41535, n41534, n38986, n41628, n41627, n41630, n41402, 
        n41413, n41537, n41409, n41508, n41509, n41510, n41308, 
        n41536;
    
    LUT4 i21062_2_lut (.A(size_d[1]), .B(sign_extend_d), .Z(n23666)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i21062_2_lut.init = 16'h6666;
    LUT4 instruction_31__I_0_188_i9_2_lut_rep_428 (.A(\instruction_d[30] ), 
         .B(\instruction_d[31] ), .Z(n41515)) /* synthesis lut_function=(A+!(B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(383[20:71])
    defparam instruction_31__I_0_188_i9_2_lut_rep_428.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_376_3_lut (.A(\instruction_d[30] ), .B(\instruction_d[31] ), 
         .C(\logic_op_d[3] ), .Z(n41463)) /* synthesis lut_function=(A+!(B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(383[20:71])
    defparam i1_2_lut_rep_376_3_lut.init = 16'hbfbf;
    LUT4 i37999_2_lut_2_lut_3_lut_4_lut (.A(\instruction_d[30] ), .B(\instruction_d[31] ), 
         .C(n41499), .D(\logic_op_d[3] ), .Z(x_result_sel_csr_d)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(383[20:71])
    defparam i37999_2_lut_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i29088_2_lut_4_lut (.A(n41427), .B(n41533), .C(\logic_op_d[3] ), 
         .D(\instruction_d[0] ), .Z(n1792)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i29088_2_lut_4_lut.init = 16'hef00;
    LUT4 i29561_2_lut_4_lut (.A(n41427), .B(n41533), .C(\logic_op_d[3] ), 
         .D(\instruction_d[15] ), .Z(n1777)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i29561_2_lut_4_lut.init = 16'hef00;
    LUT4 i1_4_lut (.A(n41397), .B(n41437), .C(n41436), .D(n41434), .Z(bra)) /* synthesis lut_function=(!(A (B+!(C+!(D))))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(405[14:54])
    defparam i1_4_lut.init = 16'h7577;
    LUT4 i29611_2_lut_4_lut (.A(n41427), .B(n41533), .C(\logic_op_d[3] ), 
         .D(\instruction_d[7] ), .Z(n1785)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i29611_2_lut_4_lut.init = 16'hef00;
    LUT4 i29612_2_lut_4_lut (.A(n41427), .B(n41533), .C(\logic_op_d[3] ), 
         .D(\instruction_d[6] ), .Z(n1786)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i29612_2_lut_4_lut.init = 16'hef00;
    LUT4 i29619_2_lut_4_lut (.A(n41427), .B(n41533), .C(\logic_op_d[3] ), 
         .D(\instruction_d[5] ), .Z(n1787)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i29619_2_lut_4_lut.init = 16'hef00;
    LUT4 i29620_2_lut_4_lut (.A(n41427), .B(n41533), .C(\logic_op_d[3] ), 
         .D(\instruction_d[4] ), .Z(n1788)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i29620_2_lut_4_lut.init = 16'hef00;
    LUT4 i29627_2_lut_4_lut (.A(n41427), .B(n41533), .C(\logic_op_d[3] ), 
         .D(\instruction_d[3] ), .Z(n1789)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i29627_2_lut_4_lut.init = 16'hef00;
    LUT4 i29628_2_lut_4_lut (.A(n41427), .B(n41533), .C(\logic_op_d[3] ), 
         .D(\instruction_d[2] ), .Z(n1790)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i29628_2_lut_4_lut.init = 16'hef00;
    LUT4 i29639_2_lut_4_lut (.A(n41427), .B(n41533), .C(\logic_op_d[3] ), 
         .D(\instruction_d[1] ), .Z(n1791)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C+!(D)))) */ ;
    defparam i29639_2_lut_4_lut.init = 16'hef00;
    LUT4 instruction_30__I_0_i6_2_lut_rep_440 (.A(size_d[0]), .B(size_d[1]), 
         .Z(n41527)) /* synthesis lut_function=(A+!(B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(397[20:65])
    defparam instruction_30__I_0_i6_2_lut_rep_440.init = 16'hbbbb;
    LUT4 i36563_2_lut_3_lut (.A(size_d[0]), .B(size_d[1]), .C(\instruction_d[30] ), 
         .Z(n39110)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(397[20:65])
    defparam i36563_2_lut_3_lut.init = 16'hfbfb;
    LUT4 i29132_2_lut_rep_441 (.A(size_d[0]), .B(size_d[1]), .Z(n41528)) /* synthesis lut_function=(A (B)) */ ;
    defparam i29132_2_lut_rep_441.init = 16'h8888;
    LUT4 i29796_2_lut_rep_377_3_lut (.A(size_d[0]), .B(size_d[1]), .C(sign_extend_d), 
         .Z(n41464)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i29796_2_lut_rep_377_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_352_3_lut (.A(size_d[0]), .B(size_d[1]), .C(sign_extend_d), 
         .Z(n41439)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam i1_2_lut_rep_352_3_lut.init = 16'hf7f7;
    LUT4 i1_2_lut_3_lut (.A(size_d[0]), .B(size_d[1]), .C(sign_extend_d), 
         .Z(n39002)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(384[20:71])
    defparam i1_2_lut_3_lut.init = 16'hfbfb;
    LUT4 i38007_3_lut_4_lut_then_3_lut (.A(\instruction_d[30] ), .B(n41499), 
         .C(\instruction_d[31] ), .Z(n41538)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(393[20:68])
    defparam i38007_3_lut_4_lut_then_3_lut.init = 16'h0101;
    LUT4 i1_2_lut_rep_373_3_lut (.A(size_d[0]), .B(size_d[1]), .C(sign_extend_d), 
         .Z(n41460)) /* synthesis lut_function=(A+!(B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(384[20:71])
    defparam i1_2_lut_rep_373_3_lut.init = 16'hbfbf;
    LUT4 i29038_2_lut_rep_340_3_lut_4_lut_4_lut_3_lut (.A(size_d[0]), .B(size_d[1]), 
         .C(sign_extend_d), .Z(n41427)) /* synthesis lut_function=(A+!(B (C)+!B !(C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(384[20:71])
    defparam i29038_2_lut_rep_340_3_lut_4_lut_4_lut_3_lut.init = 16'hbebe;
    LUT4 i2_4_lut_rep_289_4_lut (.A(n41419), .B(n39002), .C(n41434), .D(bra), 
         .Z(n41376)) /* synthesis lut_function=(A+(B (D)+!B ((D)+!C))) */ ;
    defparam i2_4_lut_rep_289_4_lut.init = 16'hffab;
    LUT4 adder_op_d_I_0_1_lut_4_lut_4_lut (.A(n41419), .B(n39002), .C(n41434), 
         .D(bra), .Z(adder_op_d_N_1339)) /* synthesis lut_function=(!(A+(B (D)+!B ((D)+!C)))) */ ;
    defparam adder_op_d_I_0_1_lut_4_lut_4_lut.init = 16'h0054;
    LUT4 i1_3_lut_rep_309_4_lut (.A(\logic_op_d[3] ), .B(n41427), .C(\instruction_d[31] ), 
         .D(\instruction_d[30] ), .Z(n41396)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_3_lut_rep_309_4_lut.init = 16'h0200;
    LUT4 i1_2_lut_rep_445 (.A(\instruction_d[30] ), .B(size_d[0]), .Z(n41532)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_rep_445.init = 16'h2222;
    LUT4 i1_2_lut_rep_359_3_lut (.A(\instruction_d[30] ), .B(size_d[0]), 
         .C(\instruction_d[31] ), .Z(n41446)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_2_lut_rep_359_3_lut.init = 16'h2020;
    LUT4 instruction_31__I_0_i9_2_lut_rep_446 (.A(\instruction_d[30] ), .B(\instruction_d[31] ), 
         .Z(n41533)) /* synthesis lut_function=((B)+!A) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(393[20:68])
    defparam instruction_31__I_0_i9_2_lut_rep_446.init = 16'hdddd;
    LUT4 instruction_31__I_0_i10_2_lut_rep_346_3_lut (.A(\instruction_d[30] ), 
         .B(\instruction_d[31] ), .C(\logic_op_d[3] ), .Z(n41433)) /* synthesis lut_function=((B+(C))+!A) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(393[20:68])
    defparam instruction_31__I_0_i10_2_lut_rep_346_3_lut.init = 16'hfdfd;
    LUT4 i3_4_lut (.A(size_d[1]), .B(size_d[0]), .C(\instruction_d[30] ), 
         .D(\logic_op_d[3] ), .Z(n8)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (((D)+!C)+!B))) */ ;
    defparam i3_4_lut.init = 16'h0048;
    LUT4 i2_3_lut_rep_258_4_lut_4_lut (.A(n41361), .B(n41364), .C(n42740), 
         .D(cycles_5__N_2495), .Z(n41345)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i2_3_lut_rep_258_4_lut_4_lut.init = 16'h4000;
    LUT4 i1_2_lut_4_lut_4_lut (.A(n41361), .B(n13), .C(w_clk_cpu_enable_958), 
         .D(n41364), .Z(n18875)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;
    defparam i1_2_lut_4_lut_4_lut.init = 16'h4000;
    LUT4 i1_4_lut_adj_175 (.A(n41515), .B(n38976), .C(n41499), .D(\logic_op_d[3] ), 
         .Z(x_result_sel_sext_N_1782)) /* synthesis lut_function=(A (B)+!A (B+!(C+!(D)))) */ ;
    defparam i1_4_lut_adj_175.init = 16'hcdcc;
    LUT4 i4_4_lut (.A(n7), .B(n40446), .C(n32034), .D(n39220), .Z(x_bypass_enable_d)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam i4_4_lut.init = 16'hefff;
    LUT4 i29049_4_lut (.A(n41499), .B(n41464), .C(n41463), .D(n41434), 
         .Z(n31609)) /* synthesis lut_function=(A ((D)+!B)+!A (B (C (D))+!B (C))) */ ;
    defparam i29049_4_lut.init = 16'hfa32;
    LUT4 i36641_4_lut (.A(n41515), .B(n41439), .C(n41499), .D(\logic_op_d[3] ), 
         .Z(n39191)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i36641_4_lut.init = 16'hfaea;
    LUT4 i1_4_lut_adj_176 (.A(n39191), .B(n58), .C(n8_adj_3651), .D(n41396), 
         .Z(m_bypass_enable_d)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;
    defparam i1_4_lut_adj_176.init = 16'hfffd;
    LUT4 i1_4_lut_adj_177 (.A(size_d[1]), .B(n23), .C(size_d[0]), .D(\instruction_d[30] ), 
         .Z(n58)) /* synthesis lut_function=(!(A+!(B+!((D)+!C)))) */ ;
    defparam i1_4_lut_adj_177.init = 16'h4454;
    LUT4 i3_4_lut_adj_178 (.A(n41312), .B(size_d[0]), .C(n39162), .D(n41494), 
         .Z(n8_adj_3651)) /* synthesis lut_function=(A+(B ((D)+!C)+!B !(C))) */ ;
    defparam i3_4_lut_adj_178.init = 16'hefaf;
    LUT4 i2_3_lut (.A(\instruction_d[30] ), .B(\logic_op_d[3] ), .C(\instruction_d[31] ), 
         .Z(n10)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(365[20:68])
    defparam i2_3_lut.init = 16'hfbfb;
    PFUMX i38107 (.BLUT(n40445), .ALUT(n40444), .C0(sign_extend_d), .Z(n40446));
    LUT4 i37926_2_lut (.A(read_idx_0_d[0]), .B(n39005), .Z(eret_d)) /* synthesis lut_function=(!(A+(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(346[20:67])
    defparam i37926_2_lut.init = 16'h1111;
    LUT4 i1_4_lut_adj_179 (.A(n20), .B(read_idx_0_d[2]), .C(n6), .D(read_idx_0_d[3]), 
         .Z(n39005)) /* synthesis lut_function=(A+!(B (C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(346[20:67])
    defparam i1_4_lut_adj_179.init = 16'hbfff;
    LUT4 i2_2_lut (.A(read_idx_0_d[1]), .B(read_idx_0_d[4]), .Z(n6)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i37932_2_lut (.A(read_idx_0_d[0]), .B(n39005), .Z(bret_d)) /* synthesis lut_function=(!((B)+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(346[20:67])
    defparam i37932_2_lut.init = 16'h2222;
    PFUMX i38583 (.BLUT(n41558), .ALUT(n41559), .C0(sign_extend_d), .Z(sign_extend_immediate));
    LUT4 bus_error_d_bdd_3_lut_4_lut (.A(n41439), .B(n41463), .C(n39005), 
         .D(bus_error_d), .Z(n41199)) /* synthesis lut_function=(A ((D)+!C)+!A (((D)+!C)+!B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(383[20:71])
    defparam bus_error_d_bdd_3_lut_4_lut.init = 16'hff1f;
    LUT4 i29477_2_lut_3_lut_3_lut_4_lut (.A(n41367), .B(n41417), .C(n22236), 
         .D(\instruction_d[12] ), .Z(n2)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(440[10] 443[53])
    defparam i29477_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i29700_2_lut_3_lut_3_lut_4_lut (.A(n41367), .B(n41417), .C(n22236), 
         .D(\instruction_d[1] ), .Z(n2_adj_3)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(440[10] 443[53])
    defparam i29700_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i29652_2_lut_3_lut_3_lut_4_lut (.A(n41367), .B(n41417), .C(n22236), 
         .D(\instruction_d[2] ), .Z(n2_adj_4)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(440[10] 443[53])
    defparam i29652_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i29565_2_lut_3_lut_3_lut_4_lut (.A(n41367), .B(n41417), .C(n22236), 
         .D(\instruction_d[3] ), .Z(n2_adj_5)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(440[10] 443[53])
    defparam i29565_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i29512_2_lut_3_lut_3_lut_4_lut (.A(n41367), .B(n41417), .C(n22236), 
         .D(\instruction_d[4] ), .Z(n2_adj_6)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(440[10] 443[53])
    defparam i29512_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i29483_2_lut_3_lut_3_lut_4_lut (.A(n41367), .B(n41417), .C(n22236), 
         .D(\instruction_d[5] ), .Z(n2_adj_7)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(440[10] 443[53])
    defparam i29483_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i29418_2_lut_3_lut_3_lut_4_lut (.A(n41367), .B(n41417), .C(n22236), 
         .D(\instruction_d[6] ), .Z(n2_adj_8)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(440[10] 443[53])
    defparam i29418_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i29354_2_lut_3_lut_3_lut_4_lut (.A(n41367), .B(n41417), .C(n22236), 
         .D(\instruction_d[7] ), .Z(n2_adj_9)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(440[10] 443[53])
    defparam i29354_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i29244_2_lut_3_lut_3_lut_4_lut (.A(n41367), .B(n41417), .C(n22236), 
         .D(\instruction_d[8] ), .Z(n2_adj_10)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(440[10] 443[53])
    defparam i29244_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i29124_2_lut_3_lut_3_lut_4_lut (.A(n41367), .B(n41417), .C(n22236), 
         .D(\instruction_d[9] ), .Z(n2_adj_11)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(440[10] 443[53])
    defparam i29124_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 i28889_2_lut_3_lut_3_lut_4_lut (.A(n41367), .B(n41417), .C(n22236), 
         .D(\instruction_d[10] ), .Z(n2_adj_12)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(440[10] 443[53])
    defparam i28889_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 bypass_data_0_31__I_0_i32_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[31]), .D(\bypass_data_0[31] ), .Z(\d_result_0[31] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i32_3_lut_4_lut.init = 16'hf780;
    LUT4 i37874_2_lut_2_lut_4_lut_then_1_lut_4_lut (.A(size_d[0]), .B(n41485), 
         .C(\logic_op_d[3] ), .D(n41477), .Z(n41631)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(345[20:71])
    defparam i37874_2_lut_2_lut_4_lut_then_1_lut_4_lut.init = 16'h1000;
    LUT4 bypass_data_0_31__I_0_i31_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[30]), .D(\bypass_data_0[30] ), .Z(\d_result_0[30] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i31_3_lut_4_lut.init = 16'hf780;
    LUT4 bypass_data_0_31__I_0_i30_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[29]), .D(\bypass_data_0[29] ), .Z(\d_result_0[29] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i30_3_lut_4_lut.init = 16'hf780;
    LUT4 bypass_data_0_31__I_0_i29_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[28]), .D(\bypass_data_0[28] ), .Z(\d_result_0[28] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i29_3_lut_4_lut.init = 16'hf780;
    LUT4 bypass_data_0_31__I_0_i28_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[27]), .D(\bypass_data_0[27] ), .Z(\d_result_0[27] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i28_3_lut_4_lut.init = 16'hf780;
    LUT4 i29482_2_lut_3_lut_3_lut_4_lut (.A(n41367), .B(n41417), .C(n22236), 
         .D(\instruction_d[0] ), .Z(n2_adj_13)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(440[10] 443[53])
    defparam i29482_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 bypass_data_0_31__I_0_i27_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[26]), .D(\bypass_data_0[26] ), .Z(\d_result_0[26] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i27_3_lut_4_lut.init = 16'hf780;
    LUT4 bypass_data_0_31__I_0_i26_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[25]), .D(\bypass_data_0[25] ), .Z(\d_result_0[25] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i26_3_lut_4_lut.init = 16'hf780;
    LUT4 bypass_data_0_31__I_0_i25_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[24]), .D(\bypass_data_0[24] ), .Z(\d_result_0[24] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i25_3_lut_4_lut.init = 16'hf780;
    LUT4 bypass_data_0_31__I_0_i24_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[23]), .D(\bypass_data_0[23] ), .Z(\d_result_0[23] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i24_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_3_lut_4_lut (.A(\instruction_d[31] ), .B(n41532), .C(n23666), 
         .D(\logic_op_d[3] ), .Z(n22224)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h0008;
    LUT4 i29634_2_lut_3_lut_3_lut_4_lut (.A(n41367), .B(n41417), .C(n22236), 
         .D(\instruction_d[11] ), .Z(n2_adj_14)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(440[10] 443[53])
    defparam i29634_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 bypass_data_0_31__I_0_i23_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[22]), .D(\bypass_data_0[22] ), .Z(\d_result_0[22] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i23_3_lut_4_lut.init = 16'hf780;
    LUT4 bypass_data_0_31__I_0_i22_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[21]), .D(\bypass_data_0[21] ), .Z(\d_result_0[21] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i22_3_lut_4_lut.init = 16'hf780;
    LUT4 bypass_data_0_31__I_0_i21_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[20]), .D(\bypass_data_0[20] ), .Z(\d_result_0[20] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i21_3_lut_4_lut.init = 16'hf780;
    LUT4 bypass_data_0_31__I_0_i20_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[19]), .D(\bypass_data_0[19] ), .Z(\d_result_0[19] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i20_3_lut_4_lut.init = 16'hf780;
    LUT4 bypass_data_0_31__I_0_i19_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[18]), .D(\bypass_data_0[18] ), .Z(\d_result_0[18] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i19_3_lut_4_lut.init = 16'hf780;
    LUT4 bypass_data_0_31__I_0_i18_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[17]), .D(\bypass_data_0[17] ), .Z(\d_result_0[17] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i18_3_lut_4_lut.init = 16'hf780;
    LUT4 bypass_data_0_31__I_0_i17_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[16]), .D(\bypass_data_0[16] ), .Z(\d_result_0[16] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i17_3_lut_4_lut.init = 16'hf780;
    LUT4 bypass_data_0_31__I_0_i16_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[15]), .D(\bypass_data_0[15] ), .Z(\d_result_0[15] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i16_3_lut_4_lut.init = 16'hf780;
    LUT4 bypass_data_0_31__I_0_i15_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[14]), .D(\bypass_data_0[14] ), .Z(\d_result_0[14] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i15_3_lut_4_lut.init = 16'hf780;
    LUT4 bypass_data_0_31__I_0_i14_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[13]), .D(\bypass_data_0[13] ), .Z(\d_result_0[13] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i14_3_lut_4_lut.init = 16'hf780;
    LUT4 bypass_data_0_31__I_0_i13_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[12]), .D(\bypass_data_0[12] ), .Z(\d_result_0[12] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i13_3_lut_4_lut.init = 16'hf780;
    LUT4 bypass_data_0_31__I_0_i12_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[11]), .D(\bypass_data_0[11] ), .Z(\d_result_0[11] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i12_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_3_lut_4_lut_4_lut (.A(size_d[1]), .B(sign_extend_d), .C(n10), 
         .Z(n39042)) /* synthesis lut_function=((B+(C))+!A) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(403[25:76])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hfdfd;
    LUT4 bypass_data_0_31__I_0_i11_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[10]), .D(\bypass_data_0[10] ), .Z(\d_result_0[10] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i11_3_lut_4_lut.init = 16'hf780;
    LUT4 bypass_data_0_31__I_0_i10_3_lut_4_lut (.A(n41486), .B(n41446), 
         .C(pc_f[9]), .D(\bypass_data_0[9] ), .Z(\d_result_0[9] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i10_3_lut_4_lut.init = 16'hf780;
    LUT4 i1_2_lut_rep_447 (.A(size_d[0]), .B(n41485), .C(\logic_op_d[3] ), 
         .D(n41477), .Z(n42722)) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(345[20:71])
    defparam i1_2_lut_rep_447.init = 16'hefff;
    LUT4 bypass_data_0_31__I_0_i9_3_lut_4_lut (.A(n41486), .B(n41446), .C(pc_f[8]), 
         .D(\bypass_data_0[8] ), .Z(\d_result_0[8] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i9_3_lut_4_lut.init = 16'hf780;
    LUT4 bypass_data_0_31__I_0_i8_3_lut_4_lut (.A(n41486), .B(n41446), .C(pc_f[7]), 
         .D(\bypass_data_0[7] ), .Z(\d_result_0[7] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i8_3_lut_4_lut.init = 16'hf780;
    LUT4 bypass_data_0_31__I_0_i7_3_lut_4_lut (.A(n41486), .B(n41446), .C(pc_f[6]), 
         .D(\bypass_data_0[6] ), .Z(\d_result_0[6] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i7_3_lut_4_lut.init = 16'hf780;
    LUT4 i38011_4_lut_rep_297 (.A(n40091), .B(n41437), .C(n39042), .D(n41433), 
         .Z(n41384)) /* synthesis lut_function=(A+!(B (C)+!B (C (D)))) */ ;
    defparam i38011_4_lut_rep_297.init = 16'hafbf;
    LUT4 bypass_data_0_31__I_0_i6_3_lut_4_lut (.A(n41486), .B(n41446), .C(pc_f[5]), 
         .D(\bypass_data_0[5] ), .Z(\d_result_0[5] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i6_3_lut_4_lut.init = 16'hf780;
    LUT4 bypass_data_0_31__I_0_i5_3_lut_4_lut (.A(n41486), .B(n41446), .C(pc_f[4]), 
         .D(\bypass_data_0[4] ), .Z(\d_result_0[4] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i5_3_lut_4_lut.init = 16'hf780;
    LUT4 i29197_2_lut_3_lut_3_lut_4_lut (.A(n41367), .B(n41417), .C(n22236), 
         .D(\instruction_d[15] ), .Z(n2_adj_15)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(440[10] 443[53])
    defparam i29197_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 bypass_data_0_31__I_0_i4_3_lut_4_lut (.A(n41486), .B(n41446), .C(pc_f[3]), 
         .D(\bypass_data_0[3] ), .Z(\d_result_0[3] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i4_3_lut_4_lut.init = 16'hf780;
    LUT4 i29224_2_lut_3_lut_3_lut_4_lut (.A(n41367), .B(n41417), .C(n22236), 
         .D(\instruction_d[14] ), .Z(n2_adj_16)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(440[10] 443[53])
    defparam i29224_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    LUT4 bypass_data_0_31__I_0_i3_3_lut_4_lut (.A(n41486), .B(n41446), .C(pc_f[2]), 
         .D(\bypass_data_0[2] ), .Z(\d_result_0[2] )) /* synthesis lut_function=(A (B (C)+!B (D))+!A (D)) */ ;
    defparam bypass_data_0_31__I_0_i3_3_lut_4_lut.init = 16'hf780;
    LUT4 i29398_2_lut_3_lut_3_lut_4_lut (.A(n41367), .B(n41417), .C(n22236), 
         .D(\instruction_d[13] ), .Z(n2_adj_17)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(440[10] 443[53])
    defparam i29398_2_lut_3_lut_3_lut_4_lut.init = 16'h0d00;
    PFUMX i38438 (.BLUT(n41138), .ALUT(n41137), .C0(\instruction_d[30] ), 
          .Z(n41139));
    LUT4 mux_681_i28_3_lut_4_lut_4_lut (.A(n41407), .B(\instruction_d[11] ), 
         .C(\instruction_d[15] ), .D(sign_extend_immediate), .Z(n1765)) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam mux_681_i28_3_lut_4_lut_4_lut.init = 16'he444;
    LUT4 mux_681_i31_3_lut_4_lut_4_lut (.A(n41407), .B(\instruction_d[14] ), 
         .C(\instruction_d[15] ), .D(sign_extend_immediate), .Z(n1762)) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam mux_681_i31_3_lut_4_lut_4_lut.init = 16'he444;
    LUT4 mux_681_i30_3_lut_4_lut_4_lut (.A(n41407), .B(\instruction_d[13] ), 
         .C(\instruction_d[15] ), .D(sign_extend_immediate), .Z(n1763)) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam mux_681_i30_3_lut_4_lut_4_lut.init = 16'he444;
    LUT4 mux_681_i27_3_lut_4_lut_4_lut (.A(n41407), .B(\instruction_d[10] ), 
         .C(\instruction_d[15] ), .D(sign_extend_immediate), .Z(n1766)) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam mux_681_i27_3_lut_4_lut_4_lut.init = 16'he444;
    LUT4 mux_681_i26_3_lut_4_lut_4_lut (.A(n41407), .B(\instruction_d[9] ), 
         .C(\instruction_d[15] ), .D(sign_extend_immediate), .Z(n1767)) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam mux_681_i26_3_lut_4_lut_4_lut.init = 16'he444;
    LUT4 i38539_then_4_lut (.A(size_d[1]), .B(\instruction_d[30] ), .C(\logic_op_d[3] ), 
         .D(\instruction_d[31] ), .Z(n41535)) /* synthesis lut_function=(A (B (C))+!A !(B (C+!(D)))) */ ;
    defparam i38539_then_4_lut.init = 16'h9591;
    LUT4 mux_681_i25_3_lut_4_lut_4_lut (.A(n41407), .B(\instruction_d[8] ), 
         .C(\instruction_d[15] ), .D(sign_extend_immediate), .Z(n1768)) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam mux_681_i25_3_lut_4_lut_4_lut.init = 16'he444;
    LUT4 mux_681_i24_3_lut_4_lut_4_lut (.A(n41407), .B(\instruction_d[7] ), 
         .C(\instruction_d[15] ), .D(sign_extend_immediate), .Z(n1769)) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam mux_681_i24_3_lut_4_lut_4_lut.init = 16'he444;
    LUT4 mux_681_i23_3_lut_4_lut_4_lut (.A(n41407), .B(\instruction_d[6] ), 
         .C(\instruction_d[15] ), .D(sign_extend_immediate), .Z(n1770)) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam mux_681_i23_3_lut_4_lut_4_lut.init = 16'he444;
    LUT4 mux_681_i22_3_lut_4_lut_4_lut (.A(n41407), .B(\instruction_d[5] ), 
         .C(\instruction_d[15] ), .D(sign_extend_immediate), .Z(n1771)) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam mux_681_i22_3_lut_4_lut_4_lut.init = 16'he444;
    LUT4 mux_681_i21_3_lut_4_lut_4_lut (.A(n41407), .B(\instruction_d[4] ), 
         .C(\instruction_d[15] ), .D(sign_extend_immediate), .Z(n1772)) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam mux_681_i21_3_lut_4_lut_4_lut.init = 16'he444;
    LUT4 i29083_2_lut_rep_407 (.A(\logic_op_d[3] ), .B(\instruction_d[30] ), 
         .Z(n41494)) /* synthesis lut_function=(A (B)) */ ;
    defparam i29083_2_lut_rep_407.init = 16'h8888;
    LUT4 i37910_2_lut_rep_332_3_lut (.A(\logic_op_d[3] ), .B(\instruction_d[30] ), 
         .C(n41427), .Z(n41419)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i37910_2_lut_rep_332_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_adj_180 (.A(\logic_op_d[3] ), .B(\instruction_d[30] ), 
         .C(sign_extend_d), .Z(n23)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_180.init = 16'h8080;
    LUT4 mux_681_i20_3_lut_4_lut_4_lut (.A(n41407), .B(\instruction_d[3] ), 
         .C(\instruction_d[15] ), .D(sign_extend_immediate), .Z(n1773)) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam mux_681_i20_3_lut_4_lut_4_lut.init = 16'he444;
    LUT4 i38539_else_4_lut (.A(size_d[1]), .B(\instruction_d[30] ), .C(\logic_op_d[3] ), 
         .D(\instruction_d[31] ), .Z(n41534)) /* synthesis lut_function=(A (B (C+(D)))+!A !(B)) */ ;
    defparam i38539_else_4_lut.init = 16'h9991;
    LUT4 mux_681_i19_3_lut_4_lut_4_lut (.A(n41407), .B(\instruction_d[2] ), 
         .C(\instruction_d[15] ), .D(sign_extend_immediate), .Z(n1774)) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam mux_681_i19_3_lut_4_lut_4_lut.init = 16'he444;
    LUT4 mux_681_i18_3_lut_4_lut_4_lut (.A(n41407), .B(\instruction_d[1] ), 
         .C(\instruction_d[15] ), .D(sign_extend_immediate), .Z(n1775)) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam mux_681_i18_3_lut_4_lut_4_lut.init = 16'he444;
    LUT4 mux_681_i17_3_lut_4_lut_4_lut (.A(n41407), .B(\instruction_d[0] ), 
         .C(\instruction_d[15] ), .D(sign_extend_immediate), .Z(n1776)) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam mux_681_i17_3_lut_4_lut_4_lut.init = 16'he444;
    LUT4 mux_681_i29_3_lut_4_lut_4_lut (.A(n41407), .B(\instruction_d[12] ), 
         .C(\instruction_d[15] ), .D(sign_extend_immediate), .Z(n1764)) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;
    defparam mux_681_i29_3_lut_4_lut_4_lut.init = 16'he444;
    LUT4 instruction_15__I_0_i2_3_lut (.A(read_idx_1_d[1]), .B(\instruction_d[12] ), 
         .C(\instruction_d[31] ), .Z(\write_idx_4__N_1770[1] )) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(549[23] 551[45])
    defparam instruction_15__I_0_i2_3_lut.init = 16'hcaca;
    LUT4 i29051_2_lut_rep_280 (.A(\instruction_d[31] ), .B(bra), .Z(n41367)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i29051_2_lut_rep_280.init = 16'heeee;
    LUT4 sign_extend_d_bdd_4_lut (.A(sign_extend_d), .B(size_d[1]), .C(size_d[0]), 
         .D(n41433), .Z(n41397)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A (B (D)+!B ((D)+!C))) */ ;
    defparam sign_extend_d_bdd_4_lut.init = 16'hff09;
    LUT4 i29042_2_lut_rep_277_3_lut_4_lut_4_lut (.A(\instruction_d[31] ), 
         .B(n41532), .C(bra), .D(n41486), .Z(n41364)) /* synthesis lut_function=(!(A (B (D))+!A !(C))) */ ;
    defparam i29042_2_lut_rep_277_3_lut_4_lut_4_lut.init = 16'h72fa;
    LUT4 i1_3_lut_rep_412 (.A(size_d[0]), .B(size_d[1]), .C(sign_extend_d), 
         .Z(n41499)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(383[20:71])
    defparam i1_3_lut_rep_412.init = 16'hefef;
    LUT4 i29328_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[19]), 
         .D(n41417), .Z(n1)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29328_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29329_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[18]), 
         .D(n41417), .Z(n1_adj_18)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29329_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i1_2_lut (.A(size_d[1]), .B(size_d[0]), .Z(n38986)) /* synthesis lut_function=(A+!(B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(403[25:76])
    defparam i1_2_lut.init = 16'hbbbb;
    LUT4 i29340_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[11]), 
         .D(n41417), .Z(n1_adj_19)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29340_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i28945_3_lut_rep_307_4_lut (.A(n41437), .B(n41436), .C(n41397), 
         .D(\instruction_d[15] ), .Z(n41394)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B+!(C+!(D))))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(355[20:71])
    defparam i28945_3_lut_rep_307_4_lut.init = 16'h4f44;
    LUT4 i29351_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[1]), 
         .D(n41417), .Z(n1_adj_20)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29351_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29349_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[2]), 
         .D(n41417), .Z(n1_adj_21)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29349_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29330_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[17]), 
         .D(n41417), .Z(n1_adj_22)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29330_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i28943_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[0]), 
         .D(n41417), .Z(n1_adj_23)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i28943_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29325_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[22]), 
         .D(n41417), .Z(n1_adj_24)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29325_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29342_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[9]), 
         .D(n41417), .Z(n1_adj_25)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29342_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i38003_2_lut_rep_274_3_lut_3_lut_4_lut_2_lut (.A(\instruction_d[31] ), 
         .B(bra), .Z(n41361)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i38003_2_lut_rep_274_3_lut_3_lut_4_lut_2_lut.init = 16'h1111;
    LUT4 i29326_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[21]), 
         .D(n41417), .Z(n1_adj_26)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29326_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29347_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[4]), 
         .D(n41417), .Z(n1_adj_27)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29347_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29314_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[26]), 
         .D(n41417), .Z(n1_adj_28)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29314_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29327_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[20]), 
         .D(n41417), .Z(n1_adj_29)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29327_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i1_4_lut_then_4_lut (.A(sign_extend_d), .B(size_d[0]), .C(\logic_op_d[3] ), 
         .D(\instruction_d[30] ), .Z(n41628)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'h0080;
    LUT4 size_d_0__bdd_3_lut_4_lut (.A(n41437), .B(n41460), .C(\logic_op_d[3] ), 
         .D(\instruction_d[31] ), .Z(n41137)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;
    defparam size_d_0__bdd_3_lut_4_lut.init = 16'h0070;
    LUT4 i2_3_lut_rep_320_4_lut (.A(n41437), .B(n41460), .C(\logic_op_d[3] ), 
         .D(n41533), .Z(n41407)) /* synthesis lut_function=(A (B+((D)+!C))+!A ((D)+!C)) */ ;
    defparam i2_3_lut_rep_320_4_lut.init = 16'hff8f;
    LUT4 i29343_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[8]), 
         .D(n41417), .Z(n1_adj_30)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29343_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29348_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[3]), 
         .D(n41417), .Z(n1_adj_31)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29348_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29341_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[10]), 
         .D(n41417), .Z(n1_adj_32)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29341_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29324_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[23]), 
         .D(n41417), .Z(n1_adj_33)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29324_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i37988_3_lut_3_lut_4_lut (.A(n41437), .B(n41460), .C(n41477), 
         .D(n41397), .Z(branch_d)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A !(C+!(D)))) */ ;
    defparam i37988_3_lut_3_lut_4_lut.init = 16'h70ff;
    LUT4 i1_4_lut_else_4_lut (.A(sign_extend_d), .B(size_d[0]), .C(\logic_op_d[3] ), 
         .D(\instruction_d[30] ), .Z(n41627)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B+(C+(D))))) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'h0009;
    LUT4 i29310_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[30]), 
         .D(n41417), .Z(n1_adj_34)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29310_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29346_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[5]), 
         .D(n41417), .Z(n1_adj_35)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29346_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29312_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[28]), 
         .D(n41417), .Z(n1_adj_36)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29312_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29339_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[12]), 
         .D(n41417), .Z(n1_adj_37)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29339_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29333_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[16]), 
         .D(n41417), .Z(n1_adj_38)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29333_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29322_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[25]), 
         .D(n41417), .Z(n1_adj_39)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29322_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29335_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[14]), 
         .D(n41417), .Z(n1_adj_40)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29335_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29344_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[7]), 
         .D(n41417), .Z(n1_adj_41)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29344_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i37874_2_lut_2_lut_4_lut_else_1_lut (.A(sign_extend_d), .B(size_d[1]), 
         .C(size_d[0]), .D(n42722), .Z(n41630)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B+(C+!(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(403[25:76])
    defparam i37874_2_lut_2_lut_4_lut_else_1_lut.init = 16'hf6ff;
    LUT4 i29338_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[13]), 
         .D(n41417), .Z(n1_adj_42)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29338_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29313_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[27]), 
         .D(n41417), .Z(n1_adj_43)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29313_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 size_d_0__bdd_4_lut_38713 (.A(size_d[0]), .B(sign_extend_d), .C(size_d[1]), 
         .D(\logic_op_d[3] ), .Z(n41138)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A !(B (C)+!B !(C+!(D))))) */ ;
    defparam size_d_0__bdd_4_lut_38713.init = 16'h4340;
    LUT4 i29334_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[15]), 
         .D(n41417), .Z(n1_adj_44)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29334_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i38034_4_lut_4_lut (.A(n41466), .B(n41139), .C(n31609), .D(n32034), 
         .Z(x_result_sel_add_N_1785)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i38034_4_lut_4_lut.init = 16'h1000;
    LUT4 i29323_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[24]), 
         .D(n41417), .Z(n1_adj_45)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29323_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29345_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[6]), 
         .D(n41417), .Z(n1_adj_46)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29345_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29309_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[31]), 
         .D(n41417), .Z(n1_adj_47)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29309_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 i29311_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(bra), .C(bypass_data_1[29]), 
         .D(n41417), .Z(n1_adj_48)) /* synthesis lut_function=(!(A ((D)+!C)+!A (((D)+!C)+!B))) */ ;
    defparam i29311_2_lut_3_lut_4_lut.init = 16'h00e0;
    LUT4 interlock_I_48_4_lut_4_lut_4_lut (.A(n41384), .B(raw_x_1), .C(raw_x_0), 
         .D(n41402), .Z(interlock_N_1327)) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;
    defparam interlock_I_48_4_lut_4_lut_4_lut.init = 16'hf400;
    LUT4 interlock_I_50_4_lut_4_lut_4_lut (.A(n41384), .B(n41411), .C(raw_m_0), 
         .D(n41402), .Z(interlock_N_1333)) /* synthesis lut_function=(A (C (D))+!A (B (D)+!B (C (D)))) */ ;
    defparam interlock_I_50_4_lut_4_lut_4_lut.init = 16'hf400;
    LUT4 i37917_4_lut_4_lut (.A(n41406), .B(n41413), .C(store_d), .D(bra), 
         .Z(write_enable_N_1809)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(395[20:70])
    defparam i37917_4_lut_4_lut.init = 16'h0004;
    LUT4 i38007_3_lut_4_lut_else_3_lut (.A(\instruction_d[30] ), .B(n41439), 
         .C(n41460), .D(\instruction_d[31] ), .Z(n41537)) /* synthesis lut_function=(!(A (C+(D))+!A (B+(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(393[20:68])
    defparam i38007_3_lut_4_lut_else_3_lut.init = 16'h001b;
    LUT4 i2_2_lut_4_lut (.A(\instruction_d[30] ), .B(\instruction_d[31] ), 
         .C(n41409), .D(n39191), .Z(n7)) /* synthesis lut_function=(!(A (B (D)+!B !(C+!(D)))+!A (D))) */ ;
    defparam i2_2_lut_4_lut.init = 16'h20ff;
    LUT4 i3_4_lut_adj_181 (.A(n23666), .B(n41532), .C(\logic_op_d[3] ), 
         .D(\instruction_d[31] ), .Z(n22236)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i3_4_lut_adj_181.init = 16'h0040;
    LUT4 i1_4_lut_then_4_lut_adj_182 (.A(size_d[1]), .B(size_d[0]), .C(\instruction_d[30] ), 
         .D(\logic_op_d[3] ), .Z(n41559)) /* synthesis lut_function=(A (B+(C))+!A !(C (D))) */ ;
    defparam i1_4_lut_then_4_lut_adj_182.init = 16'hadfd;
    LUT4 i1_4_lut_else_4_lut_adj_183 (.A(size_d[1]), .B(size_d[0]), .C(\instruction_d[30] ), 
         .D(\logic_op_d[3] ), .Z(n41558)) /* synthesis lut_function=(A+(B (C)+!B (C+!(D)))) */ ;
    defparam i1_4_lut_else_4_lut_adj_183.init = 16'hfafb;
    LUT4 i1_2_lut_rep_421 (.A(\logic_op_d[3] ), .B(\instruction_d[30] ), 
         .Z(n41508)) /* synthesis lut_function=(A+(B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(374[20:65])
    defparam i1_2_lut_rep_421.init = 16'heeee;
    LUT4 i29473_2_lut_3_lut_4_lut (.A(\logic_op_d[3] ), .B(\instruction_d[30] ), 
         .C(n41509), .D(sign_extend_d), .Z(n32034)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(374[20:65])
    defparam i29473_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 i38014_2_lut_2_lut_3_lut_4_lut (.A(\logic_op_d[3] ), .B(\instruction_d[30] ), 
         .C(n41527), .D(sign_extend_d), .Z(w_result_sel_mul_d)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(374[20:65])
    defparam i38014_2_lut_2_lut_3_lut_4_lut.init = 16'h0001;
    LUT4 instruction_30__I_0_192_i6_2_lut_rep_422 (.A(size_d[0]), .B(size_d[1]), 
         .Z(n41509)) /* synthesis lut_function=((B)+!A) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(390[20:64])
    defparam instruction_30__I_0_192_i6_2_lut_rep_422.init = 16'hdddd;
    LUT4 instruction_30__I_0_196_i7_2_lut_rep_423 (.A(\logic_op_d[3] ), .B(\instruction_d[30] ), 
         .Z(n41510)) /* synthesis lut_function=((B)+!A) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(396[20:66])
    defparam instruction_30__I_0_196_i7_2_lut_rep_423.init = 16'hdddd;
    LUT4 size_d_1__bdd_3_lut_38440_4_lut (.A(\logic_op_d[3] ), .B(n41477), 
         .C(size_d[0]), .D(size_d[1]), .Z(n40445)) /* synthesis lut_function=(!(A+((C (D)+!C !(D))+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(346[20:67])
    defparam size_d_1__bdd_3_lut_38440_4_lut.init = 16'h0440;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\logic_op_d[3] ), .B(n41477), .C(sign_extend_d), 
         .D(n41528), .Z(n38976)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(346[20:67])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h4000;
    LUT4 i1_3_lut_4_lut_adj_184 (.A(\logic_op_d[3] ), .B(n41477), .C(n38986), 
         .D(sign_extend_d), .Z(n25722)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(346[20:67])
    defparam i1_3_lut_4_lut_adj_184.init = 16'hfffb;
    LUT4 size_d_1__bdd_3_lut_38106_4_lut (.A(\logic_op_d[3] ), .B(n41477), 
         .C(n41528), .D(n39110), .Z(n40444)) /* synthesis lut_function=(!(A (D)+!A !(B (C+!(D))+!B !(D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(346[20:67])
    defparam size_d_1__bdd_3_lut_38106_4_lut.init = 16'h40ff;
    LUT4 i1_2_lut_rep_315_3_lut_4_lut (.A(n41477), .B(\logic_op_d[3] ), 
         .C(n41460), .D(n41437), .Z(n41402)) /* synthesis lut_function=(((C (D))+!B)+!A) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(405[14:54])
    defparam i1_2_lut_rep_315_3_lut_4_lut.init = 16'hf777;
    LUT4 i1_2_lut_rep_322_3_lut_4_lut (.A(size_d[0]), .B(n41485), .C(\logic_op_d[3] ), 
         .D(n41460), .Z(n41409)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(345[20:71])
    defparam i1_2_lut_rep_322_3_lut_4_lut.init = 16'h10f0;
    LUT4 equal_19659_i20_2_lut_3_lut_4_lut (.A(size_d[0]), .B(n41485), .C(n41477), 
         .D(\logic_op_d[3] ), .Z(n20)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(345[20:71])
    defparam equal_19659_i20_2_lut_3_lut_4_lut.init = 16'hffef;
    LUT4 op_raise_I_0_2_lut_3_lut_4_lut (.A(sign_extend_d), .B(n41528), 
         .C(\instruction_d[2] ), .D(n41463), .Z(scall_d)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(392[20:69])
    defparam op_raise_I_0_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 i37923_2_lut_3_lut_4_lut (.A(sign_extend_d), .B(n41528), .C(\instruction_d[2] ), 
         .D(n41463), .Z(break_d)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(392[20:69])
    defparam i37923_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 n10_bdd_4_lut_38538 (.A(size_d[0]), .B(size_d[1]), .C(\instruction_d[30] ), 
         .D(\logic_op_d[3] ), .Z(n41308)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C)+!B))) */ ;
    defparam n10_bdd_4_lut_38538.init = 16'h0e04;
    PFUMX i38567 (.BLUT(n41534), .ALUT(n41535), .C0(size_d[0]), .Z(n41536));
    LUT4 n41311_bdd_3_lut (.A(n41536), .B(n41308), .C(sign_extend_d), 
         .Z(n41312)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n41311_bdd_3_lut.init = 16'hcaca;
    LUT4 i29181_4_lut (.A(read_idx_1_d[4]), .B(n41417), .C(\instruction_d[15] ), 
         .D(\instruction_d[31] ), .Z(\write_idx_d[4] )) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(547[20] 551[45])
    defparam i29181_4_lut.init = 16'hfcee;
    LUT4 i29194_4_lut (.A(read_idx_1_d[3]), .B(n41417), .C(\instruction_d[14] ), 
         .D(\instruction_d[31] ), .Z(\write_idx_d[3] )) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(547[20] 551[45])
    defparam i29194_4_lut.init = 16'hfcee;
    LUT4 i38009_2_lut_3_lut_4_lut (.A(\instruction_d[31] ), .B(n41508), 
         .C(n41464), .D(n41499), .Z(n40091)) /* synthesis lut_function=(!(A+(B+!(C+!(D))))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(365[20:68])
    defparam i38009_2_lut_3_lut_4_lut.init = 16'h1011;
    LUT4 i1_2_lut_rep_326_3_lut_4_lut (.A(\logic_op_d[3] ), .B(n41515), 
         .C(n41528), .D(sign_extend_d), .Z(n41413)) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(383[20:71])
    defparam i1_2_lut_rep_326_3_lut_4_lut.init = 16'hffdf;
    LUT4 i36615_2_lut_3_lut_4_lut (.A(sign_extend_d), .B(n41528), .C(n41477), 
         .D(\logic_op_d[3] ), .Z(n39162)) /* synthesis lut_function=((((D)+!C)+!B)+!A) */ ;
    defparam i36615_2_lut_3_lut_4_lut.init = 16'hff7f;
    LUT4 i36669_3_lut_4_lut (.A(size_d[1]), .B(n41510), .C(size_d[0]), 
         .D(sign_extend_d), .Z(n39220)) /* synthesis lut_function=(A+(B+!(C+!(D)))) */ ;
    defparam i36669_3_lut_4_lut.init = 16'hefee;
    LUT4 i29195_4_lut (.A(read_idx_1_d[2]), .B(n41417), .C(\instruction_d[13] ), 
         .D(\instruction_d[31] ), .Z(\write_idx_d[2] )) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(547[20] 551[45])
    defparam i29195_4_lut.init = 16'hfcee;
    LUT4 i1_2_lut_3_lut_4_lut_adj_185 (.A(\logic_op_d[3] ), .B(n41515), 
         .C(n41528), .D(sign_extend_d), .Z(n25724)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(380[20:70])
    defparam i1_2_lut_3_lut_4_lut_adj_185.init = 16'hffef;
    LUT4 i4_3_lut_rep_379 (.A(\instruction_d[31] ), .B(n8), .C(sign_extend_d), 
         .Z(n41466)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i4_3_lut_rep_379.init = 16'h0808;
    LUT4 sign_extend_immediate_I_0_2_lut_rep_293 (.A(sign_extend_immediate), 
         .B(\instruction_d[15] ), .Z(n41380)) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(591[34:73])
    defparam sign_extend_immediate_I_0_2_lut_rep_293.init = 16'h8888;
    LUT4 i29147_2_lut_rep_390 (.A(\instruction_d[30] ), .B(\instruction_d[31] ), 
         .Z(n41477)) /* synthesis lut_function=(A (B)) */ ;
    defparam i29147_2_lut_rep_390.init = 16'h8888;
    LUT4 equal_19659_i19_2_lut_rep_347_3_lut (.A(\instruction_d[30] ), .B(\instruction_d[31] ), 
         .C(\logic_op_d[3] ), .Z(n41434)) /* synthesis lut_function=(((C)+!B)+!A) */ ;
    defparam equal_19659_i19_2_lut_rep_347_3_lut.init = 16'hf7f7;
    LUT4 i37992_2_lut_rep_319_2_lut_3_lut_4_lut (.A(\instruction_d[30] ), 
         .B(\instruction_d[31] ), .C(n41499), .D(\logic_op_d[3] ), .Z(n41406)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;
    defparam i37992_2_lut_rep_319_2_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_rep_349_3_lut (.A(\instruction_d[30] ), .B(\instruction_d[31] ), 
         .C(\logic_op_d[3] ), .Z(n41436)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_349_3_lut.init = 16'h8080;
    LUT4 i29060_4_lut (.A(read_idx_1_d[0]), .B(n41417), .C(\instruction_d[11] ), 
         .D(\instruction_d[31] ), .Z(\write_idx_d[0] )) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(547[20] 551[45])
    defparam i29060_4_lut.init = 16'hfcee;
    PFUMX i38569 (.BLUT(n41537), .ALUT(n41538), .C0(\logic_op_d[3] ), 
          .Z(store_d));
    PFUMX i38631 (.BLUT(n41630), .ALUT(n41631), .C0(n41433), .Z(branch_predict_d));
    PFUMX i38629 (.BLUT(n41627), .ALUT(n41628), .C0(size_d[1]), .Z(m_result_sel_shift_d));
    LUT4 i1_2_lut_rep_398 (.A(sign_extend_d), .B(size_d[1]), .Z(n41485)) /* synthesis lut_function=(A+(B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(345[20:71])
    defparam i1_2_lut_rep_398.init = 16'heeee;
    LUT4 i1_2_lut_rep_350_3_lut (.A(sign_extend_d), .B(size_d[1]), .C(size_d[0]), 
         .Z(n41437)) /* synthesis lut_function=(A+(B+(C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_decoder.v(345[20:71])
    defparam i1_2_lut_rep_350_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_399 (.A(sign_extend_d), .B(size_d[1]), .Z(n41486)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_399.init = 16'h8888;
    LUT4 i1_2_lut_rep_330_3_lut_4_lut (.A(sign_extend_d), .B(size_d[1]), 
         .C(n41532), .D(\instruction_d[31] ), .Z(n41417)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_rep_330_3_lut_4_lut.init = 16'h8000;
    
endmodule
//
// Verilog Description of module lm32_adder
//

module lm32_adder (muliplicand, operand_1_x, adder_op_x, adder_op_x_n, 
            adder_result_x, adder_carry_n_x) /* synthesis syn_module_defined=1 */ ;
    input [31:0]muliplicand;
    input [31:0]operand_1_x;
    input adder_op_x;
    input adder_op_x_n;
    output [31:0]adder_result_x;
    output adder_carry_n_x;
    
    
    lm32_addsub addsub (.muliplicand({muliplicand}), .operand_1_x({operand_1_x}), 
            .adder_op_x(adder_op_x), .adder_op_x_n(adder_op_x_n), .adder_result_x({adder_result_x}), 
            .adder_carry_n_x(adder_carry_n_x)) /* synthesis syn_module_defined=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_adder.v(100[13] 109[6])
    
endmodule
//
// Verilog Description of module lm32_addsub
//

module lm32_addsub (muliplicand, operand_1_x, adder_op_x, adder_op_x_n, 
            adder_result_x, adder_carry_n_x) /* synthesis syn_module_defined=1 */ ;
    input [31:0]muliplicand;
    input [31:0]operand_1_x;
    input adder_op_x;
    input adder_op_x_n;
    output [31:0]adder_result_x;
    output adder_carry_n_x;
    
    
    pmi_addsubMo32324b7f59e pmi_addsubMachXO2off3232 (.DataA({muliplicand}), 
            .DataB({operand_1_x}), .Result({adder_result_x}), .Cin(adder_op_x), 
            .Add_Sub(adder_op_x_n), .Cout(adder_carry_n_x)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=20, LSE_LCOL=13, LSE_RCOL=6, LSE_LLINE=100, LSE_RLINE=109 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_adder.v(100[13] 109[6])
    defparam pmi_addsubMachXO2off3232.module_type = "pmi_addsub";
    defparam pmi_addsubMachXO2off3232.pmi_family = "MachXO2";
    defparam pmi_addsubMachXO2off3232.pmi_sign = "off";
    defparam pmi_addsubMachXO2off3232.pmi_result_width = 32;
    defparam pmi_addsubMachXO2off3232.pmi_data_width = 32;
    
endmodule
//
// Verilog Description of module lm32_monitor
//

module lm32_monitor (data, ROM_DAT_O, w_clk_cpu, n87, \counter[2] , 
            \LM32D_DAT_O[15] , \SHAREDBUS_SEL_I[1] , n41490, ROM_ACK_O, 
            n42726, \data[21] , \LM32D_DAT_O[14] , \LM32D_DAT_O[13] , 
            \LM32D_DAT_O[12] , \LM32D_DAT_O[11] , \data[19] , \LM32D_DAT_O[10] , 
            \LM32D_DAT_O[9] , w_clk_cpu_enable_303, \data[30] , \LM32D_DAT_O[8] , 
            \LM32D_DAT_O[7] , n41426, \LM32D_DAT_O[0] , \LM32D_DAT_O[6] , 
            \data[29] , \data[28] , n93, n92, n41422, n41435, n35, 
            \data[27] , \data[26] , \data[25] , \data[18] , \data[24] , 
            \LM32D_DAT_O[5] , \LM32D_DAT_O[4] , \LM32D_DAT_O[3] , \LM32D_DAT_O[2] , 
            \data[23] , \LM32D_DAT_O[1] , \data[17] , \data[16] , n96, 
            \data[22] , \data[20] , GND_net, \SHAREDBUS_ADR_I[10] , 
            \SHAREDBUS_ADR_I[9] , \SHAREDBUS_ADR_I[8] , \SHAREDBUS_ADR_I[7] , 
            \SHAREDBUS_ADR_I[6] , \SHAREDBUS_ADR_I[5] , \SHAREDBUS_ADR_I[4] , 
            \SHAREDBUS_ADR_I[3] , \SHAREDBUS_ADR_I[2] , VCC_net, counter_2__N_178) /* synthesis syn_module_defined=1 */ ;
    output [31:0]data;
    output [31:0]ROM_DAT_O;
    input w_clk_cpu;
    input [7:0]n87;
    input \counter[2] ;
    input \LM32D_DAT_O[15] ;
    input \SHAREDBUS_SEL_I[1] ;
    input n41490;
    output ROM_ACK_O;
    input n42726;
    output \data[21] ;
    input \LM32D_DAT_O[14] ;
    input \LM32D_DAT_O[13] ;
    input \LM32D_DAT_O[12] ;
    input \LM32D_DAT_O[11] ;
    output \data[19] ;
    input \LM32D_DAT_O[10] ;
    input \LM32D_DAT_O[9] ;
    input w_clk_cpu_enable_303;
    output \data[30] ;
    input \LM32D_DAT_O[8] ;
    input \LM32D_DAT_O[7] ;
    input n41426;
    input \LM32D_DAT_O[0] ;
    input \LM32D_DAT_O[6] ;
    output \data[29] ;
    output \data[28] ;
    input [0:0]n93;
    input [0:0]n92;
    output n41422;
    input n41435;
    input n35;
    output \data[27] ;
    output \data[26] ;
    output \data[25] ;
    output \data[18] ;
    output \data[24] ;
    input \LM32D_DAT_O[5] ;
    input \LM32D_DAT_O[4] ;
    input \LM32D_DAT_O[3] ;
    input \LM32D_DAT_O[2] ;
    output \data[23] ;
    input \LM32D_DAT_O[1] ;
    output \data[17] ;
    output \data[16] ;
    input [7:0]n96;
    output \data[22] ;
    output \data[20] ;
    input GND_net;
    input \SHAREDBUS_ADR_I[10] ;
    input \SHAREDBUS_ADR_I[9] ;
    input \SHAREDBUS_ADR_I[8] ;
    input \SHAREDBUS_ADR_I[7] ;
    input \SHAREDBUS_ADR_I[6] ;
    input \SHAREDBUS_ADR_I[5] ;
    input \SHAREDBUS_ADR_I[4] ;
    input \SHAREDBUS_ADR_I[3] ;
    input \SHAREDBUS_ADR_I[2] ;
    input VCC_net;
    input counter_2__N_178;
    
    wire w_clk_cpu /* synthesis SET_AS_NETWORK=w_clk_cpu, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(22[6:15])
    wire [1:0]state;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(104[11:16])
    wire [31:0]n20632;
    
    wire w_clk_cpu_enable_679, n22505;
    wire [31:0]data_c;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(105[23:27])
    wire [31:0]write_data;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(107[22:32])
    
    wire w_clk_cpu_enable_980;
    wire [7:0]n78;
    
    wire n41525, w_clk_cpu_enable_175, w_clk_cpu_enable_178, n35807;
    wire [7:0]n69;
    
    wire write_enable;
    
    LUT4 i28990_2_lut (.A(data[31]), .B(state[0]), .Z(n20632[31])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i28990_2_lut.init = 16'h8888;
    FD1P3IX MON_DAT_O__i20 (.D(n20632[20]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[20])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i20.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i2 (.D(n20632[2]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[2])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i2.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i19 (.D(n20632[19]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[19])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i19.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i1 (.D(n20632[1]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[1])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i1.GSR = "DISABLED";
    LUT4 i29022_2_lut (.A(data_c[15]), .B(state[0]), .Z(n20632[15])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29022_2_lut.init = 16'h8888;
    LUT4 i29023_2_lut (.A(data_c[14]), .B(state[0]), .Z(n20632[14])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29023_2_lut.init = 16'h8888;
    FD1P3IX MON_DAT_O__i18 (.D(n20632[18]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[18])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i18.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i17 (.D(n20632[17]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[17])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i17.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i16 (.D(n20632[16]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[16])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i16.GSR = "DISABLED";
    FD1P3AX write_data_i0_i17 (.D(n87[1]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[17])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i17.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i0 (.D(n20632[0]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[0])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i0.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i31 (.D(n20632[31]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[31])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i31.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i15 (.D(n20632[15]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[15])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i15.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i14 (.D(n20632[14]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[14])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i14.GSR = "DISABLED";
    FD1P3AX write_data_i0_i16 (.D(n87[0]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[16])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i16.GSR = "DISABLED";
    FD1P3AX write_data_i0_i15 (.D(n78[7]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[15])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i15.GSR = "DISABLED";
    LUT4 i1_2_lut_rep_438 (.A(state[0]), .B(state[1]), .Z(n41525)) /* synthesis lut_function=(!((B)+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam i1_2_lut_rep_438.init = 16'h2222;
    LUT4 i2_3_lut_4_lut_3_lut (.A(state[0]), .B(state[1]), .C(w_clk_cpu_enable_175), 
         .Z(w_clk_cpu_enable_178)) /* synthesis lut_function=(A ((C)+!B)+!A (B+(C))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam i2_3_lut_4_lut_3_lut.init = 16'hf6f6;
    FD1P3AX write_data_i0_i14 (.D(n78[6]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[14])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i14.GSR = "DISABLED";
    LUT4 i1_2_lut_3_lut (.A(state[0]), .B(state[1]), .C(\counter[2] ), 
         .Z(w_clk_cpu_enable_980)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam i1_2_lut_3_lut.init = 16'h2020;
    LUT4 i33330_1_lut_2_lut (.A(state[0]), .B(state[1]), .Z(n35807)) /* synthesis lut_function=((B)+!A) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam i33330_1_lut_2_lut.init = 16'hdddd;
    FD1P3AX write_data_i0_i13 (.D(n78[5]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[13])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i13.GSR = "DISABLED";
    FD1P3AX write_data_i0_i12 (.D(n78[4]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[12])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i12.GSR = "DISABLED";
    FD1P3AX write_data_i0_i11 (.D(n78[3]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[11])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i11.GSR = "DISABLED";
    FD1P3AX write_data_i0_i10 (.D(n78[2]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[10])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i10.GSR = "DISABLED";
    FD1P3AX write_data_i0_i9 (.D(n78[1]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[9])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i9.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i30 (.D(n20632[30]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[30])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i30.GSR = "DISABLED";
    FD1P3AX write_data_i0_i8 (.D(n78[0]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[8])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i8.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i13 (.D(n20632[13]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[13])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i13.GSR = "DISABLED";
    LUT4 i29036_2_lut (.A(data_c[1]), .B(state[0]), .Z(n20632[1])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29036_2_lut.init = 16'h8888;
    FD1P3AX write_data_i0_i7 (.D(n69[7]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[7])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i7.GSR = "DISABLED";
    LUT4 mux_7_i8_4_lut (.A(data_c[15]), .B(\LM32D_DAT_O[15] ), .C(\SHAREDBUS_SEL_I[1] ), 
         .D(n41490), .Z(n78[7])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(165[36:79])
    defparam mux_7_i8_4_lut.init = 16'h0aca;
    FD1P3AX write_data_i0_i0 (.D(n69[0]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[0])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i0.GSR = "DISABLED";
    FD1S3AX MON_ACK_O_31 (.D(n41525), .CK(w_clk_cpu), .Q(ROM_ACK_O)) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_ACK_O_31.GSR = "ENABLED";
    FD1P3IX state_i0 (.D(n42726), .SP(w_clk_cpu_enable_175), .CD(w_clk_cpu_enable_679), 
            .CK(w_clk_cpu), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam state_i0.GSR = "ENABLED";
    FD1P3IX MON_DAT_O__i12 (.D(n20632[12]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[12])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i12.GSR = "DISABLED";
    FD1P3AX state_i1 (.D(n41525), .SP(w_clk_cpu_enable_178), .CK(w_clk_cpu), 
            .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam state_i1.GSR = "ENABLED";
    FD1P3AX write_data_i0_i6 (.D(n69[6]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[6])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i6.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i29 (.D(n20632[29]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[29])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i29.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i11 (.D(n20632[11]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[11])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i11.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i28 (.D(n20632[28]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[28])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i28.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i10 (.D(n20632[10]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[10])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i10.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i27 (.D(n20632[27]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[27])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i27.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i9 (.D(n20632[9]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[9])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i9.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i26 (.D(n20632[26]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[26])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i26.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i8 (.D(n20632[8]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[8])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i8.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i25 (.D(n20632[25]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[25])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i25.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i7 (.D(n20632[7]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[7])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i7.GSR = "DISABLED";
    LUT4 i29016_2_lut (.A(\data[21] ), .B(state[0]), .Z(n20632[21])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29016_2_lut.init = 16'h8888;
    LUT4 i29034_2_lut (.A(data_c[3]), .B(state[0]), .Z(n20632[3])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29034_2_lut.init = 16'h8888;
    FD1P3IX MON_DAT_O__i24 (.D(n20632[24]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[24])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i24.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i6 (.D(n20632[6]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[6])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i6.GSR = "DISABLED";
    LUT4 mux_7_i7_4_lut (.A(data_c[14]), .B(\LM32D_DAT_O[14] ), .C(\SHAREDBUS_SEL_I[1] ), 
         .D(n41490), .Z(n78[6])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(165[36:79])
    defparam mux_7_i7_4_lut.init = 16'h0aca;
    LUT4 mux_7_i6_4_lut (.A(data_c[13]), .B(\LM32D_DAT_O[13] ), .C(\SHAREDBUS_SEL_I[1] ), 
         .D(n41490), .Z(n78[5])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(165[36:79])
    defparam mux_7_i6_4_lut.init = 16'h0aca;
    FD1P3AX write_data_i0_i5 (.D(n69[5]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[5])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i5.GSR = "DISABLED";
    FD1P3AX write_data_i0_i4 (.D(n69[4]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[4])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i4.GSR = "DISABLED";
    LUT4 mux_7_i5_4_lut (.A(data_c[12]), .B(\LM32D_DAT_O[12] ), .C(\SHAREDBUS_SEL_I[1] ), 
         .D(n41490), .Z(n78[4])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(165[36:79])
    defparam mux_7_i5_4_lut.init = 16'h0aca;
    FD1P3AX write_data_i0_i3 (.D(n69[3]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[3])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i3.GSR = "DISABLED";
    LUT4 mux_7_i4_4_lut (.A(data_c[11]), .B(\LM32D_DAT_O[11] ), .C(\SHAREDBUS_SEL_I[1] ), 
         .D(n41490), .Z(n78[3])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(165[36:79])
    defparam mux_7_i4_4_lut.init = 16'h0aca;
    FD1P3AX write_data_i0_i2 (.D(n69[2]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[2])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i2.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i23 (.D(n20632[23]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[23])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i23.GSR = "DISABLED";
    LUT4 i29018_2_lut (.A(\data[19] ), .B(state[0]), .Z(n20632[19])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29018_2_lut.init = 16'h8888;
    FD1P3IX MON_DAT_O__i5 (.D(n20632[5]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[5])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i5.GSR = "DISABLED";
    FD1P3AX write_data_i0_i1 (.D(n69[1]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[1])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i1.GSR = "DISABLED";
    LUT4 mux_7_i3_4_lut (.A(data_c[10]), .B(\LM32D_DAT_O[10] ), .C(\SHAREDBUS_SEL_I[1] ), 
         .D(n41490), .Z(n78[2])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(165[36:79])
    defparam mux_7_i3_4_lut.init = 16'h0aca;
    LUT4 mux_7_i2_4_lut (.A(data_c[9]), .B(\LM32D_DAT_O[9] ), .C(\SHAREDBUS_SEL_I[1] ), 
         .D(n41490), .Z(n78[1])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(165[36:79])
    defparam mux_7_i2_4_lut.init = 16'h0aca;
    FD1P3IX write_enable_30 (.D(n42726), .SP(w_clk_cpu_enable_303), .CD(n35807), 
            .CK(w_clk_cpu), .Q(write_enable));   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_enable_30.GSR = "ENABLED";
    LUT4 i29004_2_lut (.A(\data[30] ), .B(state[0]), .Z(n20632[30])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29004_2_lut.init = 16'h8888;
    LUT4 mux_7_i1_4_lut (.A(data_c[8]), .B(\LM32D_DAT_O[8] ), .C(\SHAREDBUS_SEL_I[1] ), 
         .D(n41490), .Z(n78[0])) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (((D)+!C)+!B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(165[36:79])
    defparam mux_7_i1_4_lut.init = 16'h0aca;
    LUT4 i29024_2_lut (.A(data_c[13]), .B(state[0]), .Z(n20632[13])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29024_2_lut.init = 16'h8888;
    LUT4 mux_6_i8_4_lut (.A(data_c[7]), .B(\LM32D_DAT_O[7] ), .C(n41426), 
         .D(n41490), .Z(n69[7])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(164[35:76])
    defparam mux_6_i8_4_lut.init = 16'ha0ac;
    LUT4 mux_6_i1_4_lut (.A(data_c[0]), .B(\LM32D_DAT_O[0] ), .C(n41426), 
         .D(n41490), .Z(n69[0])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(164[35:76])
    defparam mux_6_i1_4_lut.init = 16'ha0ac;
    LUT4 i29025_2_lut (.A(data_c[12]), .B(state[0]), .Z(n20632[12])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29025_2_lut.init = 16'h8888;
    LUT4 mux_6_i7_4_lut (.A(data_c[6]), .B(\LM32D_DAT_O[6] ), .C(n41426), 
         .D(n41490), .Z(n69[6])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(164[35:76])
    defparam mux_6_i7_4_lut.init = 16'ha0ac;
    LUT4 i29005_2_lut (.A(\data[29] ), .B(state[0]), .Z(n20632[29])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29005_2_lut.init = 16'h8888;
    LUT4 i29026_2_lut (.A(data_c[11]), .B(state[0]), .Z(n20632[11])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29026_2_lut.init = 16'h8888;
    LUT4 i29009_2_lut (.A(\data[28] ), .B(state[0]), .Z(n20632[28])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29009_2_lut.init = 16'h8888;
    LUT4 i29027_2_lut (.A(data_c[10]), .B(state[0]), .Z(n20632[10])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29027_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_335 (.A(n93[0]), .B(n92[0]), .Z(n41422)) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(183[17:61])
    defparam i1_2_lut_rep_335.init = 16'h8888;
    LUT4 i1_3_lut_4_lut (.A(n93[0]), .B(n92[0]), .C(n41435), .D(n35), 
         .Z(w_clk_cpu_enable_175)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(183[17:61])
    defparam i1_3_lut_4_lut.init = 16'h0008;
    LUT4 i29010_2_lut (.A(\data[27] ), .B(state[0]), .Z(n20632[27])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29010_2_lut.init = 16'h8888;
    LUT4 i29028_2_lut (.A(data_c[9]), .B(state[0]), .Z(n20632[9])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29028_2_lut.init = 16'h8888;
    LUT4 i29011_2_lut (.A(\data[26] ), .B(state[0]), .Z(n20632[26])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29011_2_lut.init = 16'h8888;
    LUT4 i29029_2_lut (.A(data_c[8]), .B(state[0]), .Z(n20632[8])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29029_2_lut.init = 16'h8888;
    FD1P3IX MON_DAT_O__i22 (.D(n20632[22]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[22])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i22.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i4 (.D(n20632[4]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[4])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i4.GSR = "DISABLED";
    LUT4 i29012_2_lut (.A(\data[25] ), .B(state[0]), .Z(n20632[25])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29012_2_lut.init = 16'h8888;
    LUT4 i29030_2_lut (.A(data_c[7]), .B(state[0]), .Z(n20632[7])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29030_2_lut.init = 16'h8888;
    LUT4 i29019_2_lut (.A(\data[18] ), .B(state[0]), .Z(n20632[18])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29019_2_lut.init = 16'h8888;
    LUT4 i29013_2_lut (.A(\data[24] ), .B(state[0]), .Z(n20632[24])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29013_2_lut.init = 16'h8888;
    LUT4 i29031_2_lut (.A(data_c[6]), .B(state[0]), .Z(n20632[6])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29031_2_lut.init = 16'h8888;
    FD1P3IX MON_DAT_O__i21 (.D(n20632[21]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[21])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i21.GSR = "DISABLED";
    FD1P3IX MON_DAT_O__i3 (.D(n20632[3]), .SP(w_clk_cpu_enable_679), .CD(n22505), 
            .CK(w_clk_cpu), .Q(ROM_DAT_O[3])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam MON_DAT_O__i3.GSR = "DISABLED";
    LUT4 mux_6_i6_4_lut (.A(data_c[5]), .B(\LM32D_DAT_O[5] ), .C(n41426), 
         .D(n41490), .Z(n69[5])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(164[35:76])
    defparam mux_6_i6_4_lut.init = 16'ha0ac;
    LUT4 mux_6_i5_4_lut (.A(data_c[4]), .B(\LM32D_DAT_O[4] ), .C(n41426), 
         .D(n41490), .Z(n69[4])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(164[35:76])
    defparam mux_6_i5_4_lut.init = 16'ha0ac;
    LUT4 mux_6_i4_4_lut (.A(data_c[3]), .B(\LM32D_DAT_O[3] ), .C(n41426), 
         .D(n41490), .Z(n69[3])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(164[35:76])
    defparam mux_6_i4_4_lut.init = 16'ha0ac;
    LUT4 mux_6_i3_4_lut (.A(data_c[2]), .B(\LM32D_DAT_O[2] ), .C(n41426), 
         .D(n41490), .Z(n69[2])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(164[35:76])
    defparam mux_6_i3_4_lut.init = 16'ha0ac;
    LUT4 i29014_2_lut (.A(\data[23] ), .B(state[0]), .Z(n20632[23])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29014_2_lut.init = 16'h8888;
    LUT4 i29032_2_lut (.A(data_c[5]), .B(state[0]), .Z(n20632[5])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29032_2_lut.init = 16'h8888;
    LUT4 mux_6_i2_4_lut (.A(data_c[1]), .B(\LM32D_DAT_O[1] ), .C(n41426), 
         .D(n41490), .Z(n69[1])) /* synthesis lut_function=(A (B (C+!(D))+!B (C))+!A !((C+(D))+!B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(164[35:76])
    defparam mux_6_i2_4_lut.init = 16'ha0ac;
    LUT4 i29020_2_lut (.A(\data[17] ), .B(state[0]), .Z(n20632[17])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29020_2_lut.init = 16'h8888;
    LUT4 i29021_2_lut (.A(\data[16] ), .B(state[0]), .Z(n20632[16])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29021_2_lut.init = 16'h8888;
    LUT4 i29277_2_lut (.A(data_c[0]), .B(state[0]), .Z(n20632[0])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29277_2_lut.init = 16'h8888;
    FD1P3AX write_data_i0_i31 (.D(n96[7]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[31])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i31.GSR = "DISABLED";
    FD1P3AX write_data_i0_i30 (.D(n96[6]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[30])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i30.GSR = "DISABLED";
    LUT4 i37825_2_lut_rep_388 (.A(state[0]), .B(state[1]), .Z(w_clk_cpu_enable_679)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam i37825_2_lut_rep_388.init = 16'h6666;
    LUT4 i1_2_lut_3_lut_2_lut (.A(state[0]), .B(state[1]), .Z(n22505)) /* synthesis lut_function=(!(A+!(B))) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam i1_2_lut_3_lut_2_lut.init = 16'h4444;
    FD1P3AX write_data_i0_i29 (.D(n96[5]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[29])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i29.GSR = "DISABLED";
    FD1P3AX write_data_i0_i28 (.D(n96[4]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[28])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i28.GSR = "DISABLED";
    FD1P3AX write_data_i0_i27 (.D(n96[3]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[27])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i27.GSR = "DISABLED";
    LUT4 i29015_2_lut (.A(\data[22] ), .B(state[0]), .Z(n20632[22])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29015_2_lut.init = 16'h8888;
    LUT4 i29033_2_lut (.A(data_c[4]), .B(state[0]), .Z(n20632[4])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29033_2_lut.init = 16'h8888;
    FD1P3AX write_data_i0_i26 (.D(n96[2]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[26])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i26.GSR = "DISABLED";
    LUT4 i29017_2_lut (.A(\data[20] ), .B(state[0]), .Z(n20632[20])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29017_2_lut.init = 16'h8888;
    LUT4 i29035_2_lut (.A(data_c[2]), .B(state[0]), .Z(n20632[2])) /* synthesis lut_function=(A (B)) */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(154[9] 186[16])
    defparam i29035_2_lut.init = 16'h8888;
    FD1P3AX write_data_i0_i25 (.D(n96[1]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[25])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i25.GSR = "DISABLED";
    FD1P3AX write_data_i0_i24 (.D(n96[0]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[24])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i24.GSR = "DISABLED";
    FD1P3AX write_data_i0_i23 (.D(n87[7]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[23])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i23.GSR = "DISABLED";
    FD1P3AX write_data_i0_i22 (.D(n87[6]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[22])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i22.GSR = "DISABLED";
    FD1P3AX write_data_i0_i21 (.D(n87[5]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[21])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i21.GSR = "DISABLED";
    FD1P3AX write_data_i0_i20 (.D(n87[4]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[20])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i20.GSR = "DISABLED";
    FD1P3AX write_data_i0_i19 (.D(n87[3]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[19])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i19.GSR = "DISABLED";
    FD1P3AX write_data_i0_i18 (.D(n87[2]), .SP(w_clk_cpu_enable_980), .CK(w_clk_cpu), 
            .Q(write_data[18])) /* synthesis LSE_LINE_FILE_ID=34, LSE_LCOL=17, LSE_RCOL=8, LSE_LLINE=398, LSE_RLINE=413 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(153[5] 187[8])
    defparam write_data_i0_i18.GSR = "DISABLED";
    lm32_monitor_ram ram (.write_data({write_data}), .GND_net(GND_net), 
            .\SHAREDBUS_ADR_I[10] (\SHAREDBUS_ADR_I[10] ), .\SHAREDBUS_ADR_I[9] (\SHAREDBUS_ADR_I[9] ), 
            .\SHAREDBUS_ADR_I[8] (\SHAREDBUS_ADR_I[8] ), .\SHAREDBUS_ADR_I[7] (\SHAREDBUS_ADR_I[7] ), 
            .\SHAREDBUS_ADR_I[6] (\SHAREDBUS_ADR_I[6] ), .\SHAREDBUS_ADR_I[5] (\SHAREDBUS_ADR_I[5] ), 
            .\SHAREDBUS_ADR_I[4] (\SHAREDBUS_ADR_I[4] ), .\SHAREDBUS_ADR_I[3] (\SHAREDBUS_ADR_I[3] ), 
            .\SHAREDBUS_ADR_I[2] (\SHAREDBUS_ADR_I[2] ), .w_clk_cpu(w_clk_cpu), 
            .VCC_net(VCC_net), .write_enable(write_enable), .counter_2__N_178(counter_2__N_178), 
            .data({data[31], \data[30] , \data[29] , \data[28] , \data[27] , 
            \data[26] , \data[25] , \data[24] , \data[23] , \data[22] , 
            \data[21] , \data[20] , \data[19] , \data[18] , \data[17] , 
            \data[16] , data_c[15:0]})) /* synthesis syn_module_defined=1 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(113[18] 130[6])
    
endmodule
//
// Verilog Description of module lm32_monitor_ram
//

module lm32_monitor_ram (write_data, GND_net, \SHAREDBUS_ADR_I[10] , \SHAREDBUS_ADR_I[9] , 
            \SHAREDBUS_ADR_I[8] , \SHAREDBUS_ADR_I[7] , \SHAREDBUS_ADR_I[6] , 
            \SHAREDBUS_ADR_I[5] , \SHAREDBUS_ADR_I[4] , \SHAREDBUS_ADR_I[3] , 
            \SHAREDBUS_ADR_I[2] , w_clk_cpu, VCC_net, write_enable, 
            counter_2__N_178, data) /* synthesis syn_module_defined=1 */ ;
    input [31:0]write_data;
    input GND_net;
    input \SHAREDBUS_ADR_I[10] ;
    input \SHAREDBUS_ADR_I[9] ;
    input \SHAREDBUS_ADR_I[8] ;
    input \SHAREDBUS_ADR_I[7] ;
    input \SHAREDBUS_ADR_I[6] ;
    input \SHAREDBUS_ADR_I[5] ;
    input \SHAREDBUS_ADR_I[4] ;
    input \SHAREDBUS_ADR_I[3] ;
    input \SHAREDBUS_ADR_I[2] ;
    input w_clk_cpu;
    input VCC_net;
    input write_enable;
    input counter_2__N_178;
    output [31:0]data;
    
    wire w_clk_cpu /* synthesis SET_AS_NETWORK=w_clk_cpu, is_clock=1 */ ;   // e:/projects/prj_fpga_lattice/prj_ve-lcmxo27000hc/lcmx_prj/projects/mico_cpu/vga_leds.v(22[6:15])
    
    DP8KC \genblk1.lm32_monitor_ram_0_3_0  (.DIA0(write_data[27]), .DIA1(write_data[28]), 
          .DIA2(write_data[29]), .DIA3(write_data[30]), .DIA4(write_data[31]), 
          .DIA5(GND_net), .DIA6(GND_net), .DIA7(GND_net), .DIA8(GND_net), 
          .ADA0(VCC_net), .ADA1(GND_net), .ADA2(GND_net), .ADA3(\SHAREDBUS_ADR_I[2] ), 
          .ADA4(\SHAREDBUS_ADR_I[3] ), .ADA5(\SHAREDBUS_ADR_I[4] ), .ADA6(\SHAREDBUS_ADR_I[5] ), 
          .ADA7(\SHAREDBUS_ADR_I[6] ), .ADA8(\SHAREDBUS_ADR_I[7] ), .ADA9(\SHAREDBUS_ADR_I[8] ), 
          .ADA10(\SHAREDBUS_ADR_I[9] ), .ADA11(\SHAREDBUS_ADR_I[10] ), .ADA12(GND_net), 
          .CEA(VCC_net), .OCEA(VCC_net), .CLKA(w_clk_cpu), .WEA(write_enable), 
          .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), .RSTA(counter_2__N_178), 
          .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), .DIB3(GND_net), 
          .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), .DIB7(GND_net), 
          .DIB8(GND_net), .ADB0(VCC_net), .ADB1(GND_net), .ADB2(GND_net), 
          .ADB3(GND_net), .ADB4(GND_net), .ADB5(GND_net), .ADB6(GND_net), 
          .ADB7(GND_net), .ADB8(GND_net), .ADB9(GND_net), .ADB10(GND_net), 
          .ADB11(GND_net), .ADB12(GND_net), .CEB(GND_net), .OCEB(GND_net), 
          .CLKB(w_clk_cpu), .WEB(GND_net), .CSB0(GND_net), .CSB1(GND_net), 
          .CSB2(GND_net), .RSTB(counter_2__N_178), .DOA0(data[27]), .DOA1(data[28]), 
          .DOA2(data[29]), .DOA3(data[30]), .DOA4(data[31])) /* synthesis MEM_LPC_FILE="lm32_monitor_ram.lpc", MEM_INIT_FILE="lm32_monitor.mem", syn_instantiated=1, LSE_LINE_FILE_ID=35, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=113, LSE_RLINE=130 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(113[18] 130[6])
    defparam \genblk1.lm32_monitor_ram_0_3_0 .DATA_WIDTH_A = 9;
    defparam \genblk1.lm32_monitor_ram_0_3_0 .DATA_WIDTH_B = 9;
    defparam \genblk1.lm32_monitor_ram_0_3_0 .REGMODE_A = "NOREG";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .REGMODE_B = "NOREG";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .CSDECODE_A = "0b000";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .CSDECODE_B = "0b000";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .WRITEMODE_A = "NORMAL";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .WRITEMODE_B = "NORMAL";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .GSR = "ENABLED";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .RESETMODE = "SYNC";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .ASYNC_RESET_RELEASE = "SYNC";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INIT_DATA = "STATIC";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_00 = "0x0381F00C170161F02E130381F00C170161F02E130381F00C170161F02E1300C0600C0600C1F03413";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_01 = "0x0381F00C170161F02E130381F00C170161F02E130381F00C170161F02E130381F00C170161F02E13";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_02 = "0x0160B0160B0160B0160B0160B0160B0160B0160B0160B0160B0160B0160B01613016060380600C17";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_03 = "0x00A0500A1800C170160B00A0B00000000000000400C0B0240B0240B0240B0240B0240B0160B0160B";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_04 = "0x03405034050340500A0500A0500A0500A0500A0500A0500A0500A0500A0500A0500A0500A0500A05";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_05 = "0x00A0500A0500A0500A0500A0500A0500A0500A0500A0500A0500A0500A0500A0500A1800A0503405";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_06 = "0x016060301A016120300801E1A01612008180081A010040241800A050340503405034050340500A05";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_07 = "0x0160B0160B016060300600A1F0101F0101F0101F0100B016060300600A0500C1F00C1F00C1F00C1F";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_08 = "0x00C0B01E0801E0801E0801E0801E0801E1703E0700E0F01E1A00C0B0241A00C0B024170160B0160B";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_09 = "0x02408028120381F02E0801E0801E1703E1800C0500A0500A0500A0500A0500C0600C1A00C0600C1A";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_0A = "0x03E170381A0160F0100F0100F0100F0100F0100F0100F0100F0100F0100F0100F02E1F02E1F03817";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_0B = "0x0381A0381A0381A038170241C00C0600C1F0120602E1F02E1F0380603E060100900C1703E1703E1C";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_0C = "0x000000000000000000000000000000000000001C0341C0341C0341C03E060381A0381A0381A0381A";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_3_0 .INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC \genblk1.lm32_monitor_ram_0_1_2  (.DIA0(write_data[9]), .DIA1(write_data[10]), 
          .DIA2(write_data[11]), .DIA3(write_data[12]), .DIA4(write_data[13]), 
          .DIA5(write_data[14]), .DIA6(write_data[15]), .DIA7(write_data[16]), 
          .DIA8(write_data[17]), .ADA0(VCC_net), .ADA1(GND_net), .ADA2(GND_net), 
          .ADA3(\SHAREDBUS_ADR_I[2] ), .ADA4(\SHAREDBUS_ADR_I[3] ), .ADA5(\SHAREDBUS_ADR_I[4] ), 
          .ADA6(\SHAREDBUS_ADR_I[5] ), .ADA7(\SHAREDBUS_ADR_I[6] ), .ADA8(\SHAREDBUS_ADR_I[7] ), 
          .ADA9(\SHAREDBUS_ADR_I[8] ), .ADA10(\SHAREDBUS_ADR_I[9] ), .ADA11(\SHAREDBUS_ADR_I[10] ), 
          .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(w_clk_cpu), 
          .WEA(write_enable), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
          .RSTA(counter_2__N_178), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
          .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
          .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), .ADB1(GND_net), 
          .ADB2(GND_net), .ADB3(GND_net), .ADB4(GND_net), .ADB5(GND_net), 
          .ADB6(GND_net), .ADB7(GND_net), .ADB8(GND_net), .ADB9(GND_net), 
          .ADB10(GND_net), .ADB11(GND_net), .ADB12(GND_net), .CEB(GND_net), 
          .OCEB(GND_net), .CLKB(w_clk_cpu), .WEB(GND_net), .CSB0(GND_net), 
          .CSB1(GND_net), .CSB2(GND_net), .RSTB(counter_2__N_178), .DOA0(data[9]), 
          .DOA1(data[10]), .DOA2(data[11]), .DOA3(data[12]), .DOA4(data[13]), 
          .DOA5(data[14]), .DOA6(data[15]), .DOA7(data[16]), .DOA8(data[17])) /* synthesis MEM_LPC_FILE="lm32_monitor_ram.lpc", MEM_INIT_FILE="lm32_monitor.mem", syn_instantiated=1, LSE_LINE_FILE_ID=35, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=113, LSE_RLINE=130 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(113[18] 130[6])
    defparam \genblk1.lm32_monitor_ram_0_1_2 .DATA_WIDTH_A = 9;
    defparam \genblk1.lm32_monitor_ram_0_1_2 .DATA_WIDTH_B = 9;
    defparam \genblk1.lm32_monitor_ram_0_1_2 .REGMODE_A = "NOREG";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .REGMODE_B = "NOREG";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .CSDECODE_A = "0b000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .CSDECODE_B = "0b000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .WRITEMODE_A = "NORMAL";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .WRITEMODE_B = "NORMAL";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .GSR = "ENABLED";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .RESETMODE = "SYNC";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .ASYNC_RESET_RELEASE = "SYNC";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INIT_DATA = "STATIC";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_00 = "0x00000100043000000000000001000420000000000000010004300000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_01 = "0x00000100042000000000000001000420000000000000010004200000000000000100042000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_02 = "0x10000301001000030100100003010010000301001000030100100003010010000000833FF8000670";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_03 = "0x30100100001F87000080100801008010080100801F88000880008800088000880009802000030100";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_04 = "0x20100201002010030080301001000030100100003010010000301001000030100100003010010000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_05 = "0x30100100003010010000301001000030100100003010010000301001000030100100000010020100";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_06 = "0x1007F001000FE0800000100800FE0810000100000FE8001000001802010030180301803018020080";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_07 = "0x30100100003007F00000101FF101FF101FF101FF100801007F0000010080101FF101FF101FF101FF";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_08 = "0x1007F1000010000100001000010000100083FE00300223FC801007F008801007F008441010010000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_09 = "0x0707F308383FFFF0080010000100083FE00000802008000180200800018000000000800000000080";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_0A = "0x3FE043FF800FE8000080000800008000080000800008000080000800008000080011FF059FF3FE04";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_0B = "0x3FF803FF803FF803FE04071FF00180101FF10000069FF059FF3FF803FE00100FF000343FE2C3FFFF";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_0C = "0x00000000000000000000000000000000000001FF301FF301FF301FF3FE803FF803FF803FF803FF80";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_1_2 .INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC \genblk1.lm32_monitor_ram_0_0_3  (.DIA0(write_data[0]), .DIA1(write_data[1]), 
          .DIA2(write_data[2]), .DIA3(write_data[3]), .DIA4(write_data[4]), 
          .DIA5(write_data[5]), .DIA6(write_data[6]), .DIA7(write_data[7]), 
          .DIA8(write_data[8]), .ADA0(VCC_net), .ADA1(GND_net), .ADA2(GND_net), 
          .ADA3(\SHAREDBUS_ADR_I[2] ), .ADA4(\SHAREDBUS_ADR_I[3] ), .ADA5(\SHAREDBUS_ADR_I[4] ), 
          .ADA6(\SHAREDBUS_ADR_I[5] ), .ADA7(\SHAREDBUS_ADR_I[6] ), .ADA8(\SHAREDBUS_ADR_I[7] ), 
          .ADA9(\SHAREDBUS_ADR_I[8] ), .ADA10(\SHAREDBUS_ADR_I[9] ), .ADA11(\SHAREDBUS_ADR_I[10] ), 
          .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(w_clk_cpu), 
          .WEA(write_enable), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
          .RSTA(counter_2__N_178), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
          .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
          .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), .ADB1(GND_net), 
          .ADB2(GND_net), .ADB3(GND_net), .ADB4(GND_net), .ADB5(GND_net), 
          .ADB6(GND_net), .ADB7(GND_net), .ADB8(GND_net), .ADB9(GND_net), 
          .ADB10(GND_net), .ADB11(GND_net), .ADB12(GND_net), .CEB(GND_net), 
          .OCEB(GND_net), .CLKB(w_clk_cpu), .WEB(GND_net), .CSB0(GND_net), 
          .CSB1(GND_net), .CSB2(GND_net), .RSTB(counter_2__N_178), .DOA0(data[0]), 
          .DOA1(data[1]), .DOA2(data[2]), .DOA3(data[3]), .DOA4(data[4]), 
          .DOA5(data[5]), .DOA6(data[6]), .DOA7(data[7]), .DOA8(data[8])) /* synthesis MEM_LPC_FILE="lm32_monitor_ram.lpc", MEM_INIT_FILE="lm32_monitor.mem", syn_instantiated=1, LSE_LINE_FILE_ID=35, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=113, LSE_RLINE=130 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(113[18] 130[6])
    defparam \genblk1.lm32_monitor_ram_0_0_3 .DATA_WIDTH_A = 9;
    defparam \genblk1.lm32_monitor_ram_0_0_3 .DATA_WIDTH_B = 9;
    defparam \genblk1.lm32_monitor_ram_0_0_3 .REGMODE_A = "NOREG";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .REGMODE_B = "NOREG";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .CSDECODE_A = "0b000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .CSDECODE_B = "0b000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .WRITEMODE_A = "NORMAL";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .WRITEMODE_B = "NORMAL";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .GSR = "ENABLED";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .RESETMODE = "SYNC";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .ASYNC_RESET_RELEASE = "SYNC";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INIT_DATA = "STATIC";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_00 = "0x10CDC008001082A000000CCE400800108320000012CEC008001083A0000000000000000003E00000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_01 = "0x07CBC008001080A0000008CC400800108120000009CCC008001081A000000ACD4008001082200000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_02 = "0x0D0640C05C0B0540A04C090440803C070340602C050240401C030140200C010000006038A003E800";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_03 = "0x0200C010003400000878000880020100201002FF34094000900008C0009C00098000800F8740E06C";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_04 = "0x00094000900008C100780E06C0D0640C05C0B0540A04C090440803C070340602C050240401C03014";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_05 = "0x0E06C0D0640C05C0B0540A04C090440803C070340602C050240401C030140200C010000E88400098";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_06 = "0x009F4000003FE00000020A8003FE001FE001FE003FD00000000E8840009800094000900008C0F878";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_07 = "0x0281803820049DC00008009DD011DF013E1015E301608009F80000C00808011E7013E9015EB017ED";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_08 = "0x003F30C65009A470DA460E42C0AE1F0EE003780000000000000A9FF000000A9FF000000080801810";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_09 = "0x001FB000003ADB2000040144100C0033400048040100C020140301C0402400000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_0A = "0x31A003680036C1B06C1A05E190701807013066120661106610066090660806607001890019C3F200";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_0B = "0x324003280032C0038200001FB002010015B02E0000170001723F6012D401001AB000002F6002FBB1";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_0C = "0x00000000000000000000000000000000000001810018300185001872944F314003180031C0032000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_0_3 .INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    DP8KC \genblk1.lm32_monitor_ram_0_2_1  (.DIA0(write_data[18]), .DIA1(write_data[19]), 
          .DIA2(write_data[20]), .DIA3(write_data[21]), .DIA4(write_data[22]), 
          .DIA5(write_data[23]), .DIA6(write_data[24]), .DIA7(write_data[25]), 
          .DIA8(write_data[26]), .ADA0(VCC_net), .ADA1(GND_net), .ADA2(GND_net), 
          .ADA3(\SHAREDBUS_ADR_I[2] ), .ADA4(\SHAREDBUS_ADR_I[3] ), .ADA5(\SHAREDBUS_ADR_I[4] ), 
          .ADA6(\SHAREDBUS_ADR_I[5] ), .ADA7(\SHAREDBUS_ADR_I[6] ), .ADA8(\SHAREDBUS_ADR_I[7] ), 
          .ADA9(\SHAREDBUS_ADR_I[8] ), .ADA10(\SHAREDBUS_ADR_I[9] ), .ADA11(\SHAREDBUS_ADR_I[10] ), 
          .ADA12(GND_net), .CEA(VCC_net), .OCEA(VCC_net), .CLKA(w_clk_cpu), 
          .WEA(write_enable), .CSA0(GND_net), .CSA1(GND_net), .CSA2(GND_net), 
          .RSTA(counter_2__N_178), .DIB0(GND_net), .DIB1(GND_net), .DIB2(GND_net), 
          .DIB3(GND_net), .DIB4(GND_net), .DIB5(GND_net), .DIB6(GND_net), 
          .DIB7(GND_net), .DIB8(GND_net), .ADB0(VCC_net), .ADB1(GND_net), 
          .ADB2(GND_net), .ADB3(GND_net), .ADB4(GND_net), .ADB5(GND_net), 
          .ADB6(GND_net), .ADB7(GND_net), .ADB8(GND_net), .ADB9(GND_net), 
          .ADB10(GND_net), .ADB11(GND_net), .ADB12(GND_net), .CEB(GND_net), 
          .OCEB(GND_net), .CLKB(w_clk_cpu), .WEB(GND_net), .CSB0(GND_net), 
          .CSB1(GND_net), .CSB2(GND_net), .RSTB(counter_2__N_178), .DOA0(data[18]), 
          .DOA1(data[19]), .DOA2(data[20]), .DOA3(data[21]), .DOA4(data[22]), 
          .DOA5(data[23]), .DOA6(data[24]), .DOA7(data[25]), .DOA8(data[26])) /* synthesis MEM_LPC_FILE="lm32_monitor_ram.lpc", MEM_INIT_FILE="lm32_monitor.mem", syn_instantiated=1, LSE_LINE_FILE_ID=35, LSE_LCOL=18, LSE_RCOL=6, LSE_LLINE=113, LSE_RLINE=130 */ ;   // E:/projects/prj_fpga_lattice/prj_VE-LCMXO27000HC/lcmx_prj/projects/mico_cpu/mico_cpu/soc/../components/lm32_top/rtl/verilog/lm32_monitor.v(113[18] 130[6])
    defparam \genblk1.lm32_monitor_ram_0_2_1 .DATA_WIDTH_A = 9;
    defparam \genblk1.lm32_monitor_ram_0_2_1 .DATA_WIDTH_B = 9;
    defparam \genblk1.lm32_monitor_ram_0_2_1 .REGMODE_A = "NOREG";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .REGMODE_B = "NOREG";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .CSDECODE_A = "0b000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .CSDECODE_B = "0b000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .WRITEMODE_A = "NORMAL";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .WRITEMODE_B = "NORMAL";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .GSR = "ENABLED";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .RESETMODE = "SYNC";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .ASYNC_RESET_RELEASE = "SYNC";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INIT_DATA = "STATIC";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_00 = "0x00000210E01CE001D00000000210E01CE001D00000000210E01CE001D00020100201002000001000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_01 = "0x00000210E01CE001D00000000210E01CE001D00000000210E01CE001D00000000210E01CE001D000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_02 = "0x1DCEE1DAED1DAED1D8EC1D8EC1D6EB1D6EB1D4EA1D4EA1D2E91D2E91D0E81D0001D1EF1FF073CEE8";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_03 = "0x1C0E01C0E83DEE81D0E81D0E80100801008010083D0E8000E8090E8070E8020E8010EF1DEEF1DCEE";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_04 = "0x00EE709EE707EE71CEE71CCE61CCE61CAE51CAE51C8E41C8E41C6E31C6E31C4E21C4E21C2E11C2E1";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_05 = "0x1CCE61CCE61CAE51CAE51C8E41C8E41C6E31C6E31C4E21C4E21C2E11C2E11C0E01C0F01CEE701EE7";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_06 = "0x1CFE71D070220701D1082107022070010E802078210100F0F81CEE701EE700EE709EE707EE71CEE7";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_07 = "0x1C6E31C6E31C5E71D1E71CEFF1C0FF1C0FF1C0FF1C0E01CFE71D1E71CEE01C0FF1C0FF1C0FF1C0FF";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_08 = "0x201082210822108221082210822108210081FE840F60400670201080E070201080E0081CEE41C8E4";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_09 = "0x0A10C0E6301FEFF0E10822108210081FEE83CEE71C8E41C8E31C6E31C6E220100200202010020018";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_0A = "0x1FE881FEDA2111021110211102111021110211102111021110211102111021108010FF010FF1FE70";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_0B = "0x1FE4A1FE421FE3A1FE70060FF2C75A0B0FF2C703010FF010FF1FF5A1FF630B163206081FE081FEFF";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_0C = "0x00000000000000000000000000000000000000FF1A4FF184FF134FF1FF001FECA1FE921FE8A1FE82";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    defparam \genblk1.lm32_monitor_ram_0_2_1 .INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000";
    
endmodule
//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

/* Verilog netlist generated by SCUBA Diamond (64-bit) 3.10.1.112 */
/* Module Version: 3.5 */
/* D:/dev/lattice/lscc/diamond/3.10_x64/ispfpga/bin/nt64/scuba -w -arch xo2c00 -n pmi_addsubMo32324b7f59e -bb -bus_exp 7 -type addsub -width 32 -unsigned -port ci -port co -pmi -lang verilog  */
/* Thu Nov 30 05:38:42 2017 */


`timescale 1 ns / 1 ps
module pmi_addsubMo32324b7f59e (DataA, DataB, Cin, Add_Sub, Result, Cout, 
    Overflow)/* synthesis NGD_DRC_MASK=1 */;
    input wire [31:0] DataA;
    input wire [31:0] DataB;
    input wire Cin;
    input wire Add_Sub;
    output wire [31:0] Result;
    output wire Cout;
    output wire Overflow;

    wire scuba_vhi;
    wire precin;
    wire ci_k;
    wire co0;
    wire co1;
    wire co2;
    wire co3;
    wire co4;
    wire co5;
    wire co6;
    wire co7;
    wire co8;
    wire co9;
    wire co10;
    wire co11;
    wire co12;
    wire co13;
    wire co14;
    wire co15;
    wire add_sub_inv;
    wire co16d;
    wire co16;
    wire scuba_vlo;

    VHI scuba_vhi_inst (.Z(scuba_vhi));

    XNOR2 XNOR2_t0 (.A(Cin), .B(Add_Sub), .Z(ci_k));

    INV INV_0 (.A(Add_Sub), .Z(add_sub_inv));

    FADD2B precin_inst102 (.A0(scuba_vlo), .A1(scuba_vlo), .B0(scuba_vlo), 
        .B1(scuba_vlo), .CI(scuba_vlo), .COUT(precin), .S0(), .S1());

    FADSU2 addsub_0 (.A0(Cin), .A1(DataA[0]), .B0(ci_k), .B1(DataB[0]), 
        .BCI(precin), .CON(Add_Sub), .BCO(co0), .S0(), .S1(Result[0]));

    FADSU2 addsub_1 (.A0(DataA[1]), .A1(DataA[2]), .B0(DataB[1]), .B1(DataB[2]), 
        .BCI(co0), .CON(Add_Sub), .BCO(co1), .S0(Result[1]), .S1(Result[2]));

    FADSU2 addsub_2 (.A0(DataA[3]), .A1(DataA[4]), .B0(DataB[3]), .B1(DataB[4]), 
        .BCI(co1), .CON(Add_Sub), .BCO(co2), .S0(Result[3]), .S1(Result[4]));

    FADSU2 addsub_3 (.A0(DataA[5]), .A1(DataA[6]), .B0(DataB[5]), .B1(DataB[6]), 
        .BCI(co2), .CON(Add_Sub), .BCO(co3), .S0(Result[5]), .S1(Result[6]));

    FADSU2 addsub_4 (.A0(DataA[7]), .A1(DataA[8]), .B0(DataB[7]), .B1(DataB[8]), 
        .BCI(co3), .CON(Add_Sub), .BCO(co4), .S0(Result[7]), .S1(Result[8]));

    FADSU2 addsub_5 (.A0(DataA[9]), .A1(DataA[10]), .B0(DataB[9]), .B1(DataB[10]), 
        .BCI(co4), .CON(Add_Sub), .BCO(co5), .S0(Result[9]), .S1(Result[10]));

    FADSU2 addsub_6 (.A0(DataA[11]), .A1(DataA[12]), .B0(DataB[11]), .B1(DataB[12]), 
        .BCI(co5), .CON(Add_Sub), .BCO(co6), .S0(Result[11]), .S1(Result[12]));

    FADSU2 addsub_7 (.A0(DataA[13]), .A1(DataA[14]), .B0(DataB[13]), .B1(DataB[14]), 
        .BCI(co6), .CON(Add_Sub), .BCO(co7), .S0(Result[13]), .S1(Result[14]));

    FADSU2 addsub_8 (.A0(DataA[15]), .A1(DataA[16]), .B0(DataB[15]), .B1(DataB[16]), 
        .BCI(co7), .CON(Add_Sub), .BCO(co8), .S0(Result[15]), .S1(Result[16]));

    FADSU2 addsub_9 (.A0(DataA[17]), .A1(DataA[18]), .B0(DataB[17]), .B1(DataB[18]), 
        .BCI(co8), .CON(Add_Sub), .BCO(co9), .S0(Result[17]), .S1(Result[18]));

    FADSU2 addsub_10 (.A0(DataA[19]), .A1(DataA[20]), .B0(DataB[19]), .B1(DataB[20]), 
        .BCI(co9), .CON(Add_Sub), .BCO(co10), .S0(Result[19]), .S1(Result[20]));

    FADSU2 addsub_11 (.A0(DataA[21]), .A1(DataA[22]), .B0(DataB[21]), .B1(DataB[22]), 
        .BCI(co10), .CON(Add_Sub), .BCO(co11), .S0(Result[21]), .S1(Result[22]));

    FADSU2 addsub_12 (.A0(DataA[23]), .A1(DataA[24]), .B0(DataB[23]), .B1(DataB[24]), 
        .BCI(co11), .CON(Add_Sub), .BCO(co12), .S0(Result[23]), .S1(Result[24]));

    FADSU2 addsub_13 (.A0(DataA[25]), .A1(DataA[26]), .B0(DataB[25]), .B1(DataB[26]), 
        .BCI(co12), .CON(Add_Sub), .BCO(co13), .S0(Result[25]), .S1(Result[26]));

    FADSU2 addsub_14 (.A0(DataA[27]), .A1(DataA[28]), .B0(DataB[27]), .B1(DataB[28]), 
        .BCI(co13), .CON(Add_Sub), .BCO(co14), .S0(Result[27]), .S1(Result[28]));

    FADSU2 addsub_15 (.A0(DataA[29]), .A1(DataA[30]), .B0(DataB[29]), .B1(DataB[30]), 
        .BCI(co14), .CON(Add_Sub), .BCO(co15), .S0(Result[29]), .S1(Result[30]));

    FADSU2 addsub_16 (.A0(DataA[31]), .A1(scuba_vlo), .B0(DataB[31]), .B1(add_sub_inv), 
        .BCI(co15), .CON(Add_Sub), .BCO(co16), .S0(Result[31]), .S1(Cout));

    VLO scuba_vlo_inst (.Z(scuba_vlo));

    FADD2B addsubd (.A0(scuba_vlo), .A1(scuba_vlo), .B0(scuba_vlo), .B1(scuba_vlo), 
        .CI(co16), .COUT(), .S0(co16d), .S1());



    // exemplar begin
    // exemplar end

endmodule
